# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__a2bb2oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.505000 1.415000 3.955000 1.875000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.175000 1.210000 5.675000 1.750000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.235000 1.375000 0.730000 1.625000 ;
        RECT 0.550000 1.625000 0.730000 1.920000 ;
        RECT 0.550000 1.920000 1.880000 2.120000 ;
        RECT 1.595000 1.425000 2.015000 1.655000 ;
        RECT 1.595000 1.655000 1.880000 1.920000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.910000 1.425000 1.425000 1.750000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.823200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.970000 0.605000 1.300000 1.075000 ;
        RECT 0.970000 1.075000 2.750000 1.245000 ;
        RECT 2.420000 1.805000 2.750000 2.735000 ;
        RECT 2.490000 0.285000 2.750000 1.075000 ;
        RECT 2.500000 1.245000 2.750000 1.805000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.110000  0.085000 0.405000 1.185000 ;
      RECT 0.110000  1.815000 0.380000 2.290000 ;
      RECT 0.110000  2.290000 2.250000 2.460000 ;
      RECT 0.110000  2.460000 0.370000 3.075000 ;
      RECT 0.540000  2.630000 0.870000 3.245000 ;
      RECT 0.575000  0.265000 1.820000 0.435000 ;
      RECT 0.575000  0.435000 0.800000 1.185000 ;
      RECT 1.040000  2.460000 1.240000 3.075000 ;
      RECT 1.470000  0.435000 1.820000 0.905000 ;
      RECT 1.490000  2.630000 1.820000 3.245000 ;
      RECT 1.990000  0.085000 2.320000 0.895000 ;
      RECT 2.050000  1.825000 2.250000 2.290000 ;
      RECT 2.050000  2.460000 2.250000 2.905000 ;
      RECT 2.050000  2.905000 3.180000 3.075000 ;
      RECT 2.920000  0.085000 3.785000 0.895000 ;
      RECT 2.920000  1.825000 3.180000 2.905000 ;
      RECT 3.085000  1.075000 4.995000 1.245000 ;
      RECT 3.085000  1.245000 3.335000 1.605000 ;
      RECT 3.455000  2.045000 4.615000 2.215000 ;
      RECT 3.455000  2.215000 3.715000 3.075000 ;
      RECT 3.885000  2.385000 4.215000 3.245000 ;
      RECT 3.955000  0.305000 4.145000 1.075000 ;
      RECT 4.135000  1.245000 4.305000 1.705000 ;
      RECT 4.135000  1.705000 5.005000 1.875000 ;
      RECT 4.315000  0.085000 4.645000 0.895000 ;
      RECT 4.385000  2.215000 4.615000 2.905000 ;
      RECT 4.385000  2.905000 5.505000 3.075000 ;
      RECT 4.785000  1.875000 5.005000 2.735000 ;
      RECT 4.825000  0.305000 4.995000 1.075000 ;
      RECT 5.175000  0.085000 5.505000 1.040000 ;
      RECT 5.175000  1.920000 5.505000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_lp__a2bb2oi_2
END LIBRARY
