# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__o2111ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.845000 1.185000 5.675000 1.435000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.865000 1.185000 4.675000 1.435000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 1.185000 3.695000 1.515000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.105000 1.210000 1.775000 1.375000 ;
        RECT 1.105000 1.375000 1.990000 1.545000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.210000 0.425000 1.750000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  1.646400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 1.165000 0.935000 1.755000 ;
        RECT 0.595000 1.755000 4.190000 1.855000 ;
        RECT 0.595000 1.855000 2.575000 1.925000 ;
        RECT 0.595000 1.925000 0.865000 3.075000 ;
        RECT 0.605000 0.595000 0.935000 1.165000 ;
        RECT 1.535000 1.925000 1.725000 3.075000 ;
        RECT 2.385000 1.685000 4.190000 1.755000 ;
        RECT 2.395000 1.925000 2.575000 3.075000 ;
        RECT 3.860000 1.855000 4.190000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.175000  0.255000 1.335000 0.425000 ;
      RECT 0.175000  0.425000 0.435000 1.040000 ;
      RECT 0.175000  1.925000 0.425000 3.245000 ;
      RECT 1.035000  2.095000 1.365000 3.245000 ;
      RECT 1.115000  0.425000 1.335000 0.870000 ;
      RECT 1.115000  0.870000 2.275000 1.040000 ;
      RECT 1.505000  0.255000 3.330000 0.425000 ;
      RECT 1.505000  0.425000 1.775000 0.700000 ;
      RECT 1.895000  2.095000 2.225000 3.245000 ;
      RECT 1.945000  0.595000 2.275000 0.870000 ;
      RECT 1.945000  1.040000 2.275000 1.205000 ;
      RECT 2.570000  0.775000 3.690000 0.845000 ;
      RECT 2.570000  0.845000 5.480000 1.015000 ;
      RECT 2.755000  2.025000 3.085000 3.245000 ;
      RECT 3.000000  0.425000 3.330000 0.605000 ;
      RECT 3.430000  2.025000 3.690000 2.905000 ;
      RECT 3.430000  2.905000 4.550000 3.075000 ;
      RECT 3.500000  0.255000 3.690000 0.775000 ;
      RECT 3.860000  0.085000 4.190000 0.675000 ;
      RECT 4.360000  0.255000 4.550000 0.845000 ;
      RECT 4.360000  1.605000 5.480000 1.775000 ;
      RECT 4.360000  1.775000 4.550000 2.905000 ;
      RECT 4.720000  0.085000 5.050000 0.675000 ;
      RECT 4.720000  1.945000 5.050000 3.245000 ;
      RECT 5.220000  0.255000 5.480000 0.845000 ;
      RECT 5.220000  1.775000 5.480000 3.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_lp__o2111ai_2
END LIBRARY
