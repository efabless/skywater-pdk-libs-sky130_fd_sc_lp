# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__o31ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.210000 1.285000 1.525000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455000 1.210000 2.275000 1.525000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.035000 1.425000 3.415000 1.755000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.645000 1.415000 4.715000 1.585000 ;
        RECT 4.260000 1.210000 4.715000 1.415000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.451100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.420000 1.815000 2.855000 1.925000 ;
        RECT 2.420000 1.925000 3.775000 2.120000 ;
        RECT 2.420000 2.120000 2.750000 2.735000 ;
        RECT 2.685000 1.075000 4.080000 1.245000 ;
        RECT 2.685000 1.245000 2.855000 1.815000 ;
        RECT 3.415000 2.120000 3.775000 3.075000 ;
        RECT 3.595000 1.755000 4.705000 1.925000 ;
        RECT 3.750000 0.595000 4.080000 1.075000 ;
        RECT 4.445000 1.925000 4.705000 3.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.180000  1.695000 2.230000 1.865000 ;
      RECT 0.180000  1.865000 0.510000 3.075000 ;
      RECT 0.250000  0.315000 0.510000 0.870000 ;
      RECT 0.250000  0.870000 3.580000 0.905000 ;
      RECT 0.250000  0.905000 2.515000 1.040000 ;
      RECT 0.680000  0.085000 1.010000 0.700000 ;
      RECT 0.680000  2.035000 0.870000 3.245000 ;
      RECT 1.040000  1.865000 1.370000 3.075000 ;
      RECT 1.180000  0.315000 1.410000 0.870000 ;
      RECT 1.540000  2.035000 1.730000 2.905000 ;
      RECT 1.540000  2.905000 3.180000 3.075000 ;
      RECT 1.580000  0.085000 2.175000 0.700000 ;
      RECT 1.900000  1.865000 2.230000 2.735000 ;
      RECT 2.345000  0.285000 2.650000 0.735000 ;
      RECT 2.345000  0.735000 3.580000 0.870000 ;
      RECT 2.820000  0.085000 3.150000 0.565000 ;
      RECT 2.920000  2.290000 3.180000 2.905000 ;
      RECT 3.320000  0.255000 4.510000 0.425000 ;
      RECT 3.320000  0.425000 3.580000 0.735000 ;
      RECT 3.945000  2.095000 4.275000 3.245000 ;
      RECT 4.250000  0.425000 4.510000 1.040000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_lp__o31ai_2
END LIBRARY
