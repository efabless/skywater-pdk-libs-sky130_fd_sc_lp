# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__nand3_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.210000 0.505000 1.750000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.105000 1.425000 1.600000 1.920000 ;
        RECT 1.105000 1.920000 2.745000 2.120000 ;
        RECT 2.490000 1.425000 3.050000 1.645000 ;
        RECT 2.490000 1.645000 2.745000 1.920000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.810000 1.425000 2.320000 1.750000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.293600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.595000 0.935000 1.070000 ;
        RECT 0.675000 1.070000 0.935000 2.290000 ;
        RECT 0.675000 2.290000 2.745000 2.460000 ;
        RECT 0.675000 2.460000 0.885000 3.075000 ;
        RECT 1.555000 2.460000 2.745000 2.490000 ;
        RECT 1.555000 2.490000 1.785000 3.075000 ;
        RECT 2.455000 2.490000 2.745000 3.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.175000  0.255000 1.315000 0.425000 ;
      RECT 0.175000  0.425000 0.435000 1.040000 ;
      RECT 0.175000  1.920000 0.505000 3.245000 ;
      RECT 1.055000  2.630000 1.385000 3.245000 ;
      RECT 1.105000  0.425000 1.315000 1.085000 ;
      RECT 1.105000  1.085000 3.245000 1.255000 ;
      RECT 1.485000  0.285000 1.815000 0.745000 ;
      RECT 1.485000  0.745000 2.815000 0.915000 ;
      RECT 1.955000  2.660000 2.285000 3.245000 ;
      RECT 1.985000  0.085000 2.315000 0.575000 ;
      RECT 2.485000  0.285000 2.815000 0.745000 ;
      RECT 2.915000  1.815000 3.175000 3.245000 ;
      RECT 2.985000  0.305000 3.245000 1.085000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_lp__nand3_2
END LIBRARY
