# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__dlrbn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.575000 1.210000 2.030000 1.750000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.795000 0.340000 7.065000 1.155000 ;
        RECT 6.795000 1.155000 6.965000 1.815000 ;
        RECT 6.795000 1.815000 7.055000 2.155000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.795000 0.255000 9.035000 3.075000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.915000 1.210000 6.625000 2.155000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.210000 0.470000 2.490000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.600000 0.085000 ;
      RECT 0.000000  3.245000 9.600000 3.415000 ;
      RECT 0.110000  0.085000 0.440000 1.040000 ;
      RECT 0.140000  2.660000 0.470000 3.245000 ;
      RECT 0.610000  0.700000 0.820000 1.030000 ;
      RECT 0.640000  1.030000 0.820000 1.250000 ;
      RECT 0.640000  1.250000 1.055000 1.580000 ;
      RECT 0.640000  1.580000 0.900000 2.775000 ;
      RECT 0.640000  2.775000 1.520000 3.075000 ;
      RECT 0.810000  0.280000 1.405000 0.450000 ;
      RECT 1.075000  0.450000 1.405000 1.080000 ;
      RECT 1.115000  1.775000 1.405000 2.445000 ;
      RECT 1.235000  1.080000 1.405000 1.775000 ;
      RECT 1.575000  0.085000 1.795000 1.040000 ;
      RECT 1.690000  1.920000 1.940000 3.245000 ;
      RECT 1.965000  0.700000 2.380000 1.040000 ;
      RECT 2.130000  1.920000 2.460000 2.445000 ;
      RECT 2.200000  1.040000 2.380000 1.775000 ;
      RECT 2.200000  1.775000 2.460000 1.920000 ;
      RECT 2.210000  0.255000 3.955000 0.445000 ;
      RECT 2.210000  0.445000 2.380000 0.700000 ;
      RECT 2.550000  0.615000 4.375000 0.795000 ;
      RECT 2.550000  0.795000 2.760000 1.150000 ;
      RECT 2.700000  1.425000 3.260000 1.595000 ;
      RECT 2.700000  1.595000 2.870000 2.285000 ;
      RECT 2.700000  2.285000 4.130000 2.595000 ;
      RECT 2.930000  0.965000 3.260000 1.425000 ;
      RECT 3.040000  1.775000 5.165000 1.945000 ;
      RECT 3.040000  1.945000 3.320000 2.115000 ;
      RECT 3.440000  0.965000 5.235000 1.155000 ;
      RECT 3.515000  2.115000 3.845000 2.285000 ;
      RECT 3.800000  2.595000 4.130000 3.025000 ;
      RECT 4.310000  2.115000 4.640000 3.245000 ;
      RECT 4.545000  0.085000 4.765000 0.765000 ;
      RECT 4.710000  1.325000 5.735000 1.605000 ;
      RECT 4.835000  1.945000 5.165000 2.170000 ;
      RECT 4.935000  0.455000 5.235000 0.965000 ;
      RECT 5.465000  0.280000 5.735000 1.325000 ;
      RECT 5.525000  2.665000 5.765000 3.245000 ;
      RECT 5.565000  1.605000 5.735000 2.325000 ;
      RECT 5.565000  2.325000 7.580000 2.495000 ;
      RECT 5.935000  2.495000 6.175000 3.075000 ;
      RECT 6.295000  0.085000 6.625000 1.040000 ;
      RECT 6.345000  2.665000 6.675000 3.245000 ;
      RECT 7.145000  1.405000 8.155000 1.575000 ;
      RECT 7.225000  1.575000 7.580000 2.325000 ;
      RECT 7.225000  2.665000 7.555000 3.245000 ;
      RECT 7.285000  0.085000 7.595000 1.155000 ;
      RECT 7.750000  1.755000 8.615000 1.925000 ;
      RECT 7.750000  1.925000 8.020000 2.485000 ;
      RECT 7.765000  0.885000 8.615000 1.115000 ;
      RECT 8.285000  0.085000 8.615000 0.715000 ;
      RECT 8.305000  2.105000 8.625000 3.245000 ;
      RECT 8.365000  1.115000 8.615000 1.755000 ;
      RECT 9.205000  0.085000 9.495000 1.130000 ;
      RECT 9.205000  1.815000 9.495000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
  END
END sky130_fd_sc_lp__dlrbn_2
END LIBRARY
