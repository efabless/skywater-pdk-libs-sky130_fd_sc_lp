# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__invlp_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  5.040000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.305000 1.345000 7.415000 1.675000 ;
        RECT 1.565000 1.675000 3.235000 1.780000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.499000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.550000 1.135000 1.780000 ;
        RECT 0.965000 1.005000 6.605000 1.175000 ;
        RECT 0.965000 1.175000 1.135000 1.550000 ;
        RECT 0.965000 1.780000 1.135000 1.950000 ;
        RECT 0.965000 1.950000 6.675000 2.015000 ;
        RECT 0.965000 2.015000 3.945000 2.120000 ;
        RECT 3.555000 0.595000 3.805000 1.005000 ;
        RECT 3.775000 1.845000 6.675000 1.950000 ;
        RECT 3.775000 2.120000 3.945000 2.735000 ;
        RECT 4.495000 0.595000 4.745000 1.005000 ;
        RECT 4.635000 2.015000 4.805000 2.735000 ;
        RECT 5.275000 0.595000 5.605000 1.005000 ;
        RECT 5.495000 2.015000 5.665000 2.735000 ;
        RECT 6.275000 0.595000 6.605000 1.005000 ;
        RECT 6.345000 2.015000 6.675000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.115000  0.085000 0.365000 1.125000 ;
      RECT 0.115000  1.815000 0.365000 3.245000 ;
      RECT 0.545000  0.255000 0.795000 0.665000 ;
      RECT 0.545000  0.665000 3.375000 0.835000 ;
      RECT 0.545000  0.835000 0.795000 1.125000 ;
      RECT 0.545000  1.950000 0.795000 2.290000 ;
      RECT 0.545000  2.290000 3.595000 2.460000 ;
      RECT 0.545000  2.460000 0.795000 3.075000 ;
      RECT 0.975000  0.085000 1.305000 0.495000 ;
      RECT 0.975000  2.630000 1.305000 3.245000 ;
      RECT 1.485000  0.255000 1.655000 0.665000 ;
      RECT 1.485000  2.460000 1.655000 3.075000 ;
      RECT 1.835000  0.085000 2.165000 0.495000 ;
      RECT 1.835000  2.630000 2.085000 3.245000 ;
      RECT 2.265000  2.460000 2.595000 3.075000 ;
      RECT 2.345000  0.255000 2.515000 0.665000 ;
      RECT 2.695000  0.085000 3.025000 0.495000 ;
      RECT 2.765000  2.630000 3.095000 3.245000 ;
      RECT 3.205000  0.255000 7.105000 0.425000 ;
      RECT 3.205000  0.425000 3.375000 0.665000 ;
      RECT 3.265000  2.460000 3.595000 2.905000 ;
      RECT 3.265000  2.905000 7.025000 3.075000 ;
      RECT 3.985000  0.425000 4.315000 0.835000 ;
      RECT 4.125000  2.185000 4.455000 2.905000 ;
      RECT 4.925000  0.425000 5.095000 0.835000 ;
      RECT 4.985000  2.185000 5.315000 2.905000 ;
      RECT 5.775000  0.425000 6.105000 0.835000 ;
      RECT 5.845000  2.185000 6.175000 2.905000 ;
      RECT 6.775000  0.425000 7.105000 1.125000 ;
      RECT 6.855000  1.845000 7.025000 2.905000 ;
      RECT 7.205000  1.845000 7.535000 3.245000 ;
      RECT 7.285000  0.085000 7.535000 1.125000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_lp__invlp_8
END LIBRARY
