# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__mux2_0
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.000000 1.210000 1.775000 1.645000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.645000 0.265000 2.465000 0.500000 ;
        RECT 2.065000 2.155000 2.465000 2.705000 ;
        RECT 2.295000 0.500000 2.465000 2.155000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805000 2.045000 1.330000 2.265000 ;
        RECT 1.160000 2.265000 1.330000 2.905000 ;
        RECT 1.160000 2.905000 2.805000 3.075000 ;
        RECT 2.635000 2.320000 3.385000 2.490000 ;
        RECT 2.635000 2.490000 2.805000 2.905000 ;
        RECT 2.985000 1.515000 3.385000 2.320000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.289300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.470000 0.650000 0.700000 ;
        RECT 0.085000 0.700000 0.355000 2.435000 ;
        RECT 0.085000 2.435000 0.470000 3.045000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.525000  0.870000 2.115000 1.040000 ;
      RECT 0.525000  1.040000 0.780000 1.670000 ;
      RECT 0.640000  2.435000 0.990000 3.245000 ;
      RECT 0.830000  0.085000 1.160000 0.700000 ;
      RECT 1.565000  1.815000 2.115000 1.985000 ;
      RECT 1.565000  1.985000 1.895000 2.735000 ;
      RECT 1.845000  0.670000 2.115000 0.870000 ;
      RECT 1.945000  1.040000 2.115000 1.815000 ;
      RECT 2.635000  1.175000 3.735000 1.345000 ;
      RECT 2.635000  1.345000 2.815000 1.845000 ;
      RECT 2.735000  0.085000 3.065000 0.985000 ;
      RECT 2.975000  2.660000 3.175000 3.245000 ;
      RECT 3.235000  0.795000 3.565000 1.035000 ;
      RECT 3.235000  1.035000 3.735000 1.175000 ;
      RECT 3.345000  2.660000 3.735000 2.940000 ;
      RECT 3.565000  1.345000 3.735000 2.660000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__mux2_0
END LIBRARY
