# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__sregrbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.40000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN ASYNC
    ANTENNADIFFAREA  2.708750 ;
    ANTENNAPARTIALMETALSIDEAREA  2.541000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  7.775000 1.920000  8.065000 1.965000 ;
        RECT  7.775000 1.965000 11.425000 2.105000 ;
        RECT  7.775000 2.105000  8.065000 2.150000 ;
        RECT 11.135000 1.920000 11.425000 1.965000 ;
        RECT 11.135000 2.105000 11.425000 2.150000 ;
    END
  END ASYNC
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.560000 1.125000 1.890000 1.455000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.598500 ;
    ANTENNAPARTIALMETALSIDEAREA  0.980000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 13.055000 1.180000 13.345000 1.410000 ;
        RECT 13.130000 1.410000 13.270000 1.965000 ;
        RECT 13.130000 1.965000 13.765000 2.105000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.598500 ;
    ANTENNAPARTIALMETALSIDEAREA  0.980000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 13.595000 1.225000 14.230000 1.365000 ;
        RECT 14.015000 1.920000 14.305000 2.150000 ;
        RECT 14.090000 1.365000 14.230000 1.920000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.980000 1.180000 3.300000 1.855000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.480000 1.475000 1.315000 1.635000 ;
        RECT 0.480000 1.635000 2.450000 1.805000 ;
        RECT 2.130000 1.285000 2.450000 1.635000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.870000 1.180000 4.195000 1.515000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 14.400000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 14.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.400000 0.085000 ;
      RECT  0.000000  3.245000 14.400000 3.415000 ;
      RECT  0.115000  0.085000  0.365000 0.710000 ;
      RECT  0.130000  0.890000  1.140000 1.220000 ;
      RECT  0.130000  1.220000  0.300000 1.985000 ;
      RECT  0.130000  1.985000  2.280000 2.315000 ;
      RECT  0.130000  2.315000  0.300000 2.635000 ;
      RECT  0.130000  2.635000  0.685000 3.065000 ;
      RECT  0.545000  0.265000  0.875000 0.890000 ;
      RECT  0.865000  2.635000  1.195000 3.245000 ;
      RECT  1.105000  0.085000  1.435000 0.675000 ;
      RECT  1.685000  2.495000  2.800000 2.665000 ;
      RECT  1.685000  2.665000  2.015000 3.065000 ;
      RECT  1.975000  0.265000  2.305000 0.675000 ;
      RECT  2.135000  0.675000  2.305000 0.855000 ;
      RECT  2.135000  0.855000  2.800000 1.025000 ;
      RECT  2.630000  1.025000  2.800000 2.165000 ;
      RECT  2.630000  2.165000  3.335000 2.495000 ;
      RECT  2.645000  2.845000  2.975000 3.245000 ;
      RECT  2.795000  0.085000  3.045000 0.675000 ;
      RECT  3.155000  2.675000  3.685000 2.845000 ;
      RECT  3.155000  2.845000  3.485000 3.065000 ;
      RECT  3.225000  0.265000  3.715000 0.675000 ;
      RECT  3.515000  0.675000  3.685000 2.675000 ;
      RECT  3.865000  1.695000  4.545000 1.865000 ;
      RECT  3.865000  1.865000  4.035000 3.065000 ;
      RECT  3.905000  0.265000  4.155000 0.830000 ;
      RECT  3.905000  0.830000  4.545000 1.000000 ;
      RECT  4.215000  2.045000  4.545000 3.245000 ;
      RECT  4.335000  0.085000  4.665000 0.650000 ;
      RECT  4.375000  1.000000  4.545000 1.225000 ;
      RECT  4.375000  1.225000  4.850000 1.555000 ;
      RECT  4.375000  1.555000  4.545000 1.695000 ;
      RECT  4.725000  1.735000  5.690000 1.905000 ;
      RECT  4.725000  1.905000  5.030000 3.065000 ;
      RECT  4.845000  0.265000  5.200000 1.045000 ;
      RECT  5.030000  1.045000  5.200000 1.550000 ;
      RECT  5.030000  1.550000  5.690000 1.735000 ;
      RECT  5.240000  2.085000  6.040000 2.255000 ;
      RECT  5.240000  2.255000  5.490000 2.755000 ;
      RECT  5.405000  0.440000  6.040000 1.035000 ;
      RECT  5.670000  2.435000  6.390000 2.755000 ;
      RECT  5.870000  1.035000  6.040000 2.085000 ;
      RECT  6.220000  0.575000  6.470000 1.375000 ;
      RECT  6.220000  1.375000  7.505000 1.545000 ;
      RECT  6.220000  1.545000  6.390000 2.435000 ;
      RECT  6.570000  2.295000  6.820000 3.245000 ;
      RECT  6.580000  1.785000  6.910000 1.885000 ;
      RECT  6.580000  1.885000  7.380000 2.115000 ;
      RECT  7.050000  0.085000  7.380000 1.195000 ;
      RECT  7.050000  2.115000  7.380000 2.330000 ;
      RECT  7.050000  2.330000  8.470000 2.500000 ;
      RECT  7.050000  2.500000  7.380000 2.725000 ;
      RECT  7.175000  1.545000  7.505000 1.705000 ;
      RECT  7.595000  2.680000  7.925000 3.245000 ;
      RECT  7.745000  1.375000  8.075000 1.705000 ;
      RECT  7.745000  1.705000  8.035000 2.150000 ;
      RECT  7.870000  0.575000  8.425000 1.195000 ;
      RECT  8.220000  1.885000  8.470000 2.330000 ;
      RECT  8.220000  2.500000  8.470000 2.725000 ;
      RECT  8.255000  1.195000  8.425000 1.375000 ;
      RECT  8.255000  1.375000  9.065000 1.705000 ;
      RECT  8.255000  1.705000  8.425000 1.885000 ;
      RECT  8.635000  0.085000  8.885000 1.195000 ;
      RECT  8.700000  1.885000  9.030000 3.245000 ;
      RECT  9.245000  1.375000  9.695000 1.780000 ;
      RECT  9.605000  0.435000 10.045000 0.985000 ;
      RECT  9.605000  0.985000 11.110000 1.195000 ;
      RECT  9.640000  2.025000 10.045000 2.195000 ;
      RECT  9.640000  2.195000  9.970000 2.905000 ;
      RECT  9.875000  1.195000 10.045000 2.025000 ;
      RECT 10.420000  1.765000 10.750000 2.095000 ;
      RECT 10.580000  1.455000 12.430000 1.625000 ;
      RECT 10.580000  1.625000 10.750000 1.765000 ;
      RECT 10.580000  2.095000 10.750000 2.330000 ;
      RECT 10.580000  2.330000 11.530000 2.500000 ;
      RECT 10.655000  0.085000 10.985000 0.805000 ;
      RECT 10.690000  2.680000 11.020000 3.245000 ;
      RECT 10.780000  1.195000 11.110000 1.275000 ;
      RECT 11.165000  1.805000 11.835000 2.095000 ;
      RECT 11.165000  2.095000 11.395000 2.150000 ;
      RECT 11.200000  2.500000 11.530000 3.065000 ;
      RECT 11.445000  0.265000 11.775000 1.455000 ;
      RECT 11.710000  2.275000 12.040000 3.245000 ;
      RECT 12.005000  0.085000 12.255000 0.725000 ;
      RECT 12.100000  1.625000 12.430000 1.785000 ;
      RECT 12.255000  2.235000 12.780000 2.325000 ;
      RECT 12.255000  2.325000 13.725000 2.495000 ;
      RECT 12.255000  2.495000 12.585000 2.915000 ;
      RECT 12.435000  0.265000 12.780000 0.725000 ;
      RECT 12.610000  0.725000 12.780000 2.235000 ;
      RECT 12.965000  0.265000 13.325000 2.145000 ;
      RECT 13.395000  2.675000 13.725000 3.245000 ;
      RECT 13.505000  0.085000 13.755000 1.145000 ;
      RECT 13.555000  1.325000 13.960000 1.655000 ;
      RECT 13.555000  1.655000 13.725000 2.325000 ;
      RECT 13.905000  1.835000 14.310000 3.065000 ;
      RECT 13.935000  0.265000 14.310000 1.145000 ;
      RECT 14.140000  1.145000 14.310000 1.835000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  0.470000  3.685000 0.640000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  0.470000  5.605000 0.640000 ;
      RECT  5.435000  1.580000  5.605000 1.750000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  1.950000  8.005000 2.120000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  1.580000  9.445000 1.750000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  1.950000 11.365000 2.120000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  1.210000 13.285000 1.380000 ;
      RECT 13.115000  1.210000 13.285000 1.380000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  1.950000 14.245000 2.120000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
    LAYER met1 ;
      RECT 3.455000 0.440000 3.745000 0.485000 ;
      RECT 3.455000 0.485000 5.665000 0.625000 ;
      RECT 3.455000 0.625000 3.745000 0.670000 ;
      RECT 5.375000 0.440000 5.665000 0.485000 ;
      RECT 5.375000 0.625000 5.665000 0.670000 ;
      RECT 5.375000 1.550000 5.665000 1.595000 ;
      RECT 5.375000 1.595000 9.505000 1.735000 ;
      RECT 5.375000 1.735000 5.665000 1.780000 ;
      RECT 9.215000 1.550000 9.505000 1.595000 ;
      RECT 9.215000 1.735000 9.505000 1.780000 ;
  END
END sky130_fd_sc_lp__sregrbp_1
END LIBRARY
