# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__a2111o_lp
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.175000 5.155000 1.845000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.935000 1.175000 4.265000 1.845000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365000 1.175000 3.715000 1.845000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 1.175000 1.390000 1.845000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.855000 0.530000 1.780000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.235000 0.265000 2.845000 0.645000 ;
        RECT 2.235000 0.645000 2.405000 1.920000 ;
        RECT 2.235000 1.920000 2.755000 2.180000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 0.675000 ;
      RECT 0.115000  2.025000 0.880000 2.195000 ;
      RECT 0.115000  2.195000 0.445000 3.065000 ;
      RECT 0.710000  0.265000 1.265000 0.825000 ;
      RECT 0.710000  0.825000 2.055000 0.995000 ;
      RECT 0.710000  0.995000 0.880000 2.025000 ;
      RECT 1.135000  2.025000 1.465000 2.360000 ;
      RECT 1.135000  2.360000 3.470000 2.530000 ;
      RECT 1.135000  2.530000 1.465000 3.065000 ;
      RECT 1.725000  0.085000 2.055000 0.645000 ;
      RECT 1.725000  0.995000 2.055000 1.790000 ;
      RECT 1.835000  2.710000 2.165000 3.245000 ;
      RECT 2.585000  0.825000 5.035000 0.995000 ;
      RECT 2.585000  0.995000 2.915000 1.495000 ;
      RECT 3.095000  0.265000 3.425000 0.825000 ;
      RECT 3.140000  2.025000 3.470000 2.360000 ;
      RECT 3.140000  2.530000 3.470000 3.065000 ;
      RECT 3.670000  2.025000 5.135000 2.195000 ;
      RECT 3.670000  2.195000 4.000000 3.065000 ;
      RECT 3.885000  0.085000 4.215000 0.645000 ;
      RECT 4.200000  2.375000 4.530000 3.245000 ;
      RECT 4.705000  0.265000 5.035000 0.825000 ;
      RECT 4.805000  2.195000 5.135000 3.065000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_lp__a2111o_lp
END LIBRARY
