# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__xnor3_lp
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.465000 1.515000 0.835000 1.845000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.002000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.345000 3.030000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.689000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.730000 0.975000 8.060000 1.380000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.375000 1.180000 9.965000 2.890000 ;
        RECT 9.375000 2.890000 9.705000 3.025000 ;
        RECT 9.715000 0.640000 9.965000 1.180000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.115000  0.525000  0.445000 1.165000 ;
      RECT 0.115000  1.165000  1.505000 1.335000 ;
      RECT 0.115000  1.335000  0.285000 2.025000 ;
      RECT 0.115000  2.025000  0.570000 3.065000 ;
      RECT 0.770000  2.025000  1.100000 3.245000 ;
      RECT 0.905000  0.085000  1.155000 0.985000 ;
      RECT 1.175000  1.335000  1.505000 1.835000 ;
      RECT 1.300000  2.025000  1.865000 2.245000 ;
      RECT 1.300000  2.245000  4.735000 2.415000 ;
      RECT 1.300000  2.415000  1.630000 3.065000 ;
      RECT 1.335000  0.265000  2.295000 0.435000 ;
      RECT 1.335000  0.435000  1.505000 1.165000 ;
      RECT 1.695000  0.615000  1.945000 0.985000 ;
      RECT 1.695000  0.985000  1.865000 2.025000 ;
      RECT 2.125000  0.435000  2.295000 0.995000 ;
      RECT 2.125000  0.995000  3.075000 1.165000 ;
      RECT 2.475000  0.085000  2.725000 0.815000 ;
      RECT 2.600000  2.595000  2.930000 3.245000 ;
      RECT 2.905000  0.265000  3.895000 0.435000 ;
      RECT 2.905000  0.435000  3.075000 0.995000 ;
      RECT 3.210000  1.815000  3.540000 2.065000 ;
      RECT 3.295000  0.615000  3.545000 1.245000 ;
      RECT 3.295000  1.245000  3.830000 1.575000 ;
      RECT 3.295000  1.575000  3.540000 1.815000 ;
      RECT 3.725000  0.435000  3.895000 0.895000 ;
      RECT 3.725000  0.895000  4.595000 1.065000 ;
      RECT 3.795000  2.595000  4.125000 2.895000 ;
      RECT 3.795000  2.895000  8.065000 3.065000 ;
      RECT 4.075000  0.265000  6.475000 0.435000 ;
      RECT 4.075000  0.435000  4.245000 0.715000 ;
      RECT 4.405000  1.245000  5.105000 1.415000 ;
      RECT 4.405000  1.415000  4.735000 2.245000 ;
      RECT 4.405000  2.415000  4.735000 2.715000 ;
      RECT 4.425000  0.615000  6.125000 0.785000 ;
      RECT 4.425000  0.785000  4.595000 0.895000 ;
      RECT 4.775000  0.965000  5.105000 1.245000 ;
      RECT 4.915000  1.795000  5.615000 1.965000 ;
      RECT 4.915000  1.965000  5.085000 2.895000 ;
      RECT 5.265000  2.145000  5.595000 2.155000 ;
      RECT 5.265000  2.155000  7.005000 2.325000 ;
      RECT 5.265000  2.325000  5.595000 2.715000 ;
      RECT 5.285000  0.965000  5.615000 1.795000 ;
      RECT 5.795000  0.785000  6.125000 1.965000 ;
      RECT 6.305000  0.435000  6.475000 2.155000 ;
      RECT 6.325000  2.505000  6.655000 2.895000 ;
      RECT 6.715000  0.265000  9.185000 0.435000 ;
      RECT 6.715000  0.435000  6.965000 1.645000 ;
      RECT 6.715000  1.645000  7.185000 1.975000 ;
      RECT 6.835000  2.325000  7.715000 2.495000 ;
      RECT 7.145000  0.615000  7.535000 0.995000 ;
      RECT 7.365000  0.995000  7.535000 1.975000 ;
      RECT 7.365000  1.975000  8.065000 2.145000 ;
      RECT 7.465000  2.495000  7.715000 2.685000 ;
      RECT 7.715000  0.615000  8.645000 0.795000 ;
      RECT 7.895000  2.145000  8.065000 2.895000 ;
      RECT 8.050000  1.560000  8.645000 1.795000 ;
      RECT 8.315000  1.795000  8.645000 3.025000 ;
      RECT 8.475000  0.795000  8.645000 1.560000 ;
      RECT 8.845000  0.730000  9.535000 0.900000 ;
      RECT 8.845000  0.900000  9.175000 1.100000 ;
      RECT 8.845000  1.985000  9.175000 3.245000 ;
      RECT 8.855000  0.435000  9.185000 0.550000 ;
      RECT 9.365000  0.085000  9.535000 0.730000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_lp__xnor3_lp
END LIBRARY
