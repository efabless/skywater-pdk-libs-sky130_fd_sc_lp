# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__sdfrtn_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.44000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.510000 1.070000 2.885000 1.405000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.581700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.880000 1.815000 13.345000 3.075000 ;
        RECT 13.085000 0.295000 13.345000 1.815000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAPARTIALMETALSIDEAREA  3.451000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  7.755000 1.430000  8.715000 1.745000 ;
        RECT  7.755000 1.745000  8.025000 2.180000 ;
        RECT  8.545000 1.745000  8.715000 2.635000 ;
        RECT  8.545000 2.635000  9.265000 2.805000 ;
        RECT  9.095000 2.805000  9.265000 2.905000 ;
        RECT  9.095000 2.905000 10.315000 3.075000 ;
        RECT 10.145000 1.375000 11.040000 1.965000 ;
        RECT 10.145000 1.965000 10.315000 2.905000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.950000 0.745000 1.885000 1.095000 ;
        RECT 1.640000 1.095000 1.885000 1.955000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.055000 1.055000 2.340000 1.575000 ;
        RECT 2.055000 1.575000 2.785000 1.850000 ;
        RECT 2.055000 1.850000 2.620000 2.105000 ;
    END
  END SCE
  PIN CLK_N
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.475000 1.345000 4.645000 1.750000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.440000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 13.440000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.440000 0.085000 ;
      RECT  0.000000  3.245000 13.440000 3.415000 ;
      RECT  0.110000  0.085000  0.405000 0.690000 ;
      RECT  0.110000  1.815000  0.405000 3.245000 ;
      RECT  0.575000  0.295000  0.870000 0.565000 ;
      RECT  0.575000  0.565000  0.770000 1.815000 ;
      RECT  0.575000  1.815000  0.810000 1.965000 ;
      RECT  0.575000  1.965000  1.425000 2.275000 ;
      RECT  0.575000  2.275000  2.960000 2.445000 ;
      RECT  0.575000  2.445000  0.810000 2.495000 ;
      RECT  1.105000  2.615000  3.525000 2.785000 ;
      RECT  1.105000  2.785000  1.435000 2.965000 ;
      RECT  1.350000  0.265000  3.550000 0.435000 ;
      RECT  1.350000  0.435000  1.680000 0.545000 ;
      RECT  1.955000  2.955000  2.625000 3.245000 ;
      RECT  2.255000  0.605000  2.585000 0.685000 ;
      RECT  2.255000  0.685000  6.290000 0.795000 ;
      RECT  2.255000  0.795000  4.035000 0.855000 ;
      RECT  2.790000  2.020000  3.265000 2.195000 ;
      RECT  2.790000  2.195000  2.960000 2.275000 ;
      RECT  3.095000  1.035000  3.425000 1.205000 ;
      RECT  3.095000  1.205000  3.265000 2.020000 ;
      RECT  3.195000  2.365000  4.035000 2.430000 ;
      RECT  3.195000  2.430000  6.235000 2.600000 ;
      RECT  3.195000  2.600000  3.525000 2.615000 ;
      RECT  3.195000  2.785000  3.525000 3.065000 ;
      RECT  3.220000  0.435000  3.550000 0.515000 ;
      RECT  3.460000  1.525000  3.695000 2.195000 ;
      RECT  3.755000  2.770000  4.085000 3.245000 ;
      RECT  3.865000  0.625000  6.290000 0.685000 ;
      RECT  3.865000  0.855000  4.035000 2.365000 ;
      RECT  3.875000  0.085000  4.205000 0.455000 ;
      RECT  4.320000  1.930000  5.215000 2.260000 ;
      RECT  4.385000  0.965000  5.215000 1.165000 ;
      RECT  4.945000  0.085000  5.275000 0.455000 ;
      RECT  4.945000  2.770000  5.275000 3.245000 ;
      RECT  5.045000  1.165000  5.215000 1.930000 ;
      RECT  5.395000  0.965000  5.820000 1.125000 ;
      RECT  5.395000  1.125000  6.630000 1.295000 ;
      RECT  5.395000  1.295000  5.820000 1.815000 ;
      RECT  5.395000  1.815000  6.630000 2.150000 ;
      RECT  5.395000  2.150000  6.160000 2.260000 ;
      RECT  5.915000  2.600000  6.235000 3.020000 ;
      RECT  6.040000  0.795000  6.290000 0.955000 ;
      RECT  6.405000  2.320000  7.000000 2.350000 ;
      RECT  6.405000  2.350000  8.375000 2.520000 ;
      RECT  6.405000  2.520000  6.695000 3.020000 ;
      RECT  6.460000  0.255000  7.350000 0.510000 ;
      RECT  6.460000  0.510000  6.630000 1.125000 ;
      RECT  6.800000  0.680000  7.000000 2.320000 ;
      RECT  7.155000  2.690000  7.455000 3.245000 ;
      RECT  7.180000  0.510000  7.350000 0.720000 ;
      RECT  7.180000  0.720000  9.450000 0.890000 ;
      RECT  7.215000  1.060000  9.110000 1.260000 ;
      RECT  7.215000  1.260000  7.545000 2.145000 ;
      RECT  7.625000  2.520000  8.375000 3.020000 ;
      RECT  8.120000  0.085000  8.450000 0.550000 ;
      RECT  8.195000  1.985000  8.375000 2.350000 ;
      RECT  8.585000  2.985000  8.915000 3.245000 ;
      RECT  8.940000  1.260000  9.110000 2.265000 ;
      RECT  8.940000  2.265000  9.460000 2.465000 ;
      RECT  9.195000  0.255000 10.110000 0.455000 ;
      RECT  9.195000  0.455000  9.450000 0.720000 ;
      RECT  9.280000  0.890000  9.450000 1.755000 ;
      RECT  9.280000  1.755000  9.625000 2.085000 ;
      RECT  9.620000  0.625000  9.965000 1.025000 ;
      RECT  9.620000  1.025000 11.600000 1.205000 ;
      RECT  9.620000  1.205000  9.965000 1.295000 ;
      RECT  9.630000  2.405000  9.965000 2.735000 ;
      RECT  9.795000  1.295000  9.965000 2.405000 ;
      RECT 10.495000  2.175000 11.390000 2.505000 ;
      RECT 10.540000  2.710000 10.870000 3.245000 ;
      RECT 10.560000  0.085000 10.890000 0.855000 ;
      RECT 11.080000  2.505000 11.380000 3.075000 ;
      RECT 11.220000  1.795000 11.940000 1.965000 ;
      RECT 11.220000  1.965000 11.390000 2.175000 ;
      RECT 11.340000  1.205000 11.600000 1.495000 ;
      RECT 11.465000  0.595000 11.940000 0.855000 ;
      RECT 11.550000  2.710000 11.840000 3.245000 ;
      RECT 11.770000  0.855000 11.940000 1.795000 ;
      RECT 11.810000  2.135000 12.280000 2.415000 ;
      RECT 12.110000  0.350000 12.355000 1.265000 ;
      RECT 12.110000  1.265000 12.915000 1.595000 ;
      RECT 12.110000  1.595000 12.280000 2.135000 ;
      RECT 12.370000  2.585000 12.710000 3.245000 ;
      RECT 12.450000  1.765000 12.710000 2.585000 ;
      RECT 12.525000  0.085000 12.915000 1.095000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  1.950000  3.685000 2.120000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  1.950000  8.005000 2.120000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
    LAYER met1 ;
      RECT 3.455000 1.920000 3.745000 1.965000 ;
      RECT 3.455000 1.965000 8.065000 2.105000 ;
      RECT 3.455000 2.105000 3.745000 2.150000 ;
      RECT 7.775000 1.920000 8.065000 1.965000 ;
      RECT 7.775000 2.105000 8.065000 2.150000 ;
  END
END sky130_fd_sc_lp__sdfrtn_1
END LIBRARY
