# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__o221ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.680000 1.345000 4.015000 1.695000 ;
        RECT 3.680000 1.695000 5.670000 1.875000 ;
        RECT 5.345000 1.210000 5.670000 1.695000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.220000 1.210000 5.175000 1.525000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.350000 1.425000 2.315000 1.675000 ;
        RECT 1.505000 1.675000 2.315000 1.705000 ;
        RECT 1.505000 1.705000 3.470000 1.875000 ;
        RECT 3.140000 1.345000 3.470000 1.705000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.485000 1.210000 2.835000 1.535000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.210000 0.355000 1.750000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.293600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.595000 0.865000 1.815000 ;
        RECT 0.535000 1.815000 1.180000 1.845000 ;
        RECT 0.535000 1.845000 1.335000 2.045000 ;
        RECT 0.535000 2.045000 4.785000 2.215000 ;
        RECT 0.535000 2.215000 0.795000 3.075000 ;
        RECT 2.415000 2.215000 2.745000 2.735000 ;
        RECT 4.455000 2.215000 4.785000 2.725000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.105000  0.255000 1.235000 0.425000 ;
      RECT 0.105000  0.425000 0.365000 1.040000 ;
      RECT 0.105000  1.920000 0.365000 3.245000 ;
      RECT 0.965000  2.385000 1.815000 3.245000 ;
      RECT 1.045000  0.425000 1.235000 1.085000 ;
      RECT 1.045000  1.085000 2.315000 1.255000 ;
      RECT 1.485000  0.255000 3.715000 0.425000 ;
      RECT 1.485000  0.425000 1.815000 0.915000 ;
      RECT 1.985000  0.595000 2.315000 0.870000 ;
      RECT 1.985000  0.870000 3.345000 1.040000 ;
      RECT 1.985000  1.040000 2.315000 1.085000 ;
      RECT 1.985000  2.385000 2.245000 2.905000 ;
      RECT 1.985000  2.905000 3.175000 3.075000 ;
      RECT 2.485000  0.425000 2.695000 0.700000 ;
      RECT 2.865000  0.595000 3.345000 0.870000 ;
      RECT 2.915000  2.385000 3.175000 2.905000 ;
      RECT 3.005000  1.040000 3.345000 1.145000 ;
      RECT 3.395000  2.385000 3.725000 3.245000 ;
      RECT 3.515000  0.425000 3.715000 0.870000 ;
      RECT 3.515000  0.870000 5.575000 1.040000 ;
      RECT 3.895000  0.085000 4.225000 0.700000 ;
      RECT 4.025000  2.385000 4.285000 2.895000 ;
      RECT 4.025000  2.895000 5.145000 3.075000 ;
      RECT 4.395000  0.305000 4.625000 0.870000 ;
      RECT 4.795000  0.085000 5.125000 0.700000 ;
      RECT 4.955000  2.045000 5.145000 2.895000 ;
      RECT 5.295000  0.305000 5.575000 0.870000 ;
      RECT 5.315000  2.045000 5.645000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_lp__o221ai_2
END LIBRARY
