# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__dfsbp_lp
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.92000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.110000 0.550000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.215000 1.850000 13.805000 2.890000 ;
        RECT 13.475000 0.265000 13.805000 0.725000 ;
        RECT 13.635000 0.725000 13.805000 1.850000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.335000 0.265000 11.665000 0.725000 ;
        RECT 11.495000 0.725000 11.665000 1.180000 ;
        RECT 11.495000 1.180000 11.925000 1.780000 ;
        RECT 11.595000 1.780000 11.925000 3.020000 ;
    END
  END Q_N
  PIN SET_B
    ANTENNAGATEAREA  0.626000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 6.335000 1.920000 6.625000 1.965000 ;
        RECT 6.335000 1.965000 9.985000 2.105000 ;
        RECT 6.335000 2.105000 6.625000 2.150000 ;
        RECT 9.695000 1.920000 9.985000 1.965000 ;
        RECT 9.695000 2.105000 9.985000 2.150000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.560000 1.450000 1.890000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.920000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 13.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.920000 0.085000 ;
      RECT  0.000000  3.245000 13.920000 3.415000 ;
      RECT  0.095000  0.085000  0.425000 0.725000 ;
      RECT  0.170000  2.025000  0.500000 3.245000 ;
      RECT  0.700000  2.025000  1.030000 3.065000 ;
      RECT  0.860000  0.265000  2.090000 0.435000 ;
      RECT  0.860000  0.435000  1.215000 0.725000 ;
      RECT  0.860000  0.725000  1.030000 2.025000 ;
      RECT  1.210000  0.905000  1.740000 1.075000 ;
      RECT  1.210000  1.075000  1.380000 1.960000 ;
      RECT  1.210000  1.960000  2.460000 2.130000 ;
      RECT  1.210000  2.130000  1.625000 3.065000 ;
      RECT  1.410000  0.615000  1.740000 0.905000 ;
      RECT  1.825000  2.310000  2.155000 3.245000 ;
      RECT  1.920000  0.435000  2.090000 1.100000 ;
      RECT  1.920000  1.100000  2.810000 1.270000 ;
      RECT  2.130000  1.555000  2.460000 1.960000 ;
      RECT  2.280000  0.085000  2.450000 0.920000 ;
      RECT  2.355000  2.310000  2.685000 2.895000 ;
      RECT  2.355000  2.895000  4.545000 3.065000 ;
      RECT  2.640000  0.265000  3.840000 0.435000 ;
      RECT  2.640000  0.435000  2.810000 1.100000 ;
      RECT  2.640000  1.270000  2.810000 1.960000 ;
      RECT  2.640000  1.960000  3.335000 2.130000 ;
      RECT  2.990000  0.615000  3.320000 1.330000 ;
      RECT  2.990000  1.330000  4.520000 1.780000 ;
      RECT  3.005000  2.130000  3.335000 2.715000 ;
      RECT  3.510000  0.435000  3.840000 0.885000 ;
      RECT  3.515000  1.780000  3.685000 2.895000 ;
      RECT  3.865000  2.075000  4.870000 2.245000 ;
      RECT  3.865000  2.245000  4.195000 2.715000 ;
      RECT  4.085000  0.425000  4.335000 0.865000 ;
      RECT  4.085000  0.865000  5.515000 1.035000 ;
      RECT  4.085000  1.035000  4.870000 1.065000 ;
      RECT  4.375000  2.505000  7.585000 2.675000 ;
      RECT  4.375000  2.675000  4.545000 2.895000 ;
      RECT  4.700000  1.065000  4.870000 2.075000 ;
      RECT  4.915000  0.085000  5.165000 0.685000 ;
      RECT  4.985000  2.855000  5.315000 3.245000 ;
      RECT  5.050000  1.215000  5.865000 1.385000 ;
      RECT  5.050000  1.385000  5.380000 2.075000 ;
      RECT  5.050000  2.075000  6.215000 2.325000 ;
      RECT  5.345000  0.265000  6.470000 0.435000 ;
      RECT  5.345000  0.435000  5.515000 0.865000 ;
      RECT  5.620000  1.565000  6.215000 1.895000 ;
      RECT  5.695000  0.615000  6.120000 1.065000 ;
      RECT  5.695000  1.065000  5.865000 1.215000 ;
      RECT  6.045000  1.245000  7.205000 1.415000 ;
      RECT  6.045000  1.415000  6.215000 1.565000 ;
      RECT  6.300000  0.435000  6.470000 1.245000 ;
      RECT  6.395000  1.605000  6.665000 2.150000 ;
      RECT  6.495000  2.855000  6.825000 3.245000 ;
      RECT  6.750000  0.085000  7.080000 1.065000 ;
      RECT  6.875000  1.415000  7.205000 1.915000 ;
      RECT  7.415000  1.300000  7.745000 1.460000 ;
      RECT  7.415000  1.460000  8.580000 1.630000 ;
      RECT  7.415000  1.630000  7.585000 2.505000 ;
      RECT  7.650000  0.605000  8.095000 0.915000 ;
      RECT  7.650000  0.915000  8.930000 1.065000 ;
      RECT  7.805000  2.075000  8.135000 2.330000 ;
      RECT  7.805000  2.330000 10.140000 2.500000 ;
      RECT  7.805000  2.500000  8.135000 3.065000 ;
      RECT  7.925000  1.065000  8.930000 1.085000 ;
      RECT  8.315000  1.630000  8.580000 1.935000 ;
      RECT  8.760000  1.085000  8.930000 2.330000 ;
      RECT  8.945000  0.085000  9.275000 0.735000 ;
      RECT  9.110000  0.915000 10.615000 1.085000 ;
      RECT  9.110000  1.085000  9.375000 1.885000 ;
      RECT  9.110000  2.680000  9.440000 3.245000 ;
      RECT  9.585000  1.265000  9.955000 2.150000 ;
      RECT  9.755000  0.265000 10.085000 0.915000 ;
      RECT  9.810000  2.500000 10.140000 2.895000 ;
      RECT  9.810000  2.895000 10.965000 3.065000 ;
      RECT 10.365000  1.085000 10.615000 2.715000 ;
      RECT 10.545000  0.085000 10.875000 0.725000 ;
      RECT 10.795000  1.170000 11.125000 1.840000 ;
      RECT 10.795000  1.840000 10.965000 2.895000 ;
      RECT 11.145000  2.020000 11.395000 3.245000 ;
      RECT 11.895000  0.265000 12.275000 0.725000 ;
      RECT 12.105000  0.725000 12.275000 1.490000 ;
      RECT 12.105000  1.490000 13.320000 1.660000 ;
      RECT 12.105000  1.660000 12.485000 2.890000 ;
      RECT 12.685000  0.085000 13.015000 0.725000 ;
      RECT 12.685000  1.850000 13.015000 3.245000 ;
      RECT 12.990000  0.990000 13.320000 1.490000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  1.950000  6.565000 2.120000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  1.950000  9.925000 2.120000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
  END
END sky130_fd_sc_lp__dfsbp_lp
END LIBRARY
