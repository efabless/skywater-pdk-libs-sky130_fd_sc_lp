# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__sdfxbp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.36000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.040000 1.385000 1.850000 2.120000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.110000 1.050000 12.870000 1.220000 ;
        RECT 12.110000 1.220000 12.335000 1.875000 ;
        RECT 12.110000 1.875000 12.920000 2.205000 ;
        RECT 12.640000 0.260000 12.870000 1.050000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.555000 0.255000 14.815000 3.075000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.145000 0.755000 1.185000 ;
        RECT 0.085000 1.185000 0.805000 2.120000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.020000 0.265000 3.285000 1.485000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 7.345000 1.140000 8.550000 1.395000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 15.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 15.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 15.360000 0.085000 ;
      RECT  0.000000  3.245000 15.360000 3.415000 ;
      RECT  0.095000  0.085000  0.425000 0.975000 ;
      RECT  0.095000  2.290000  2.115000 2.460000 ;
      RECT  0.095000  2.460000  0.425000 3.075000 ;
      RECT  0.595000  2.630000  0.875000 3.245000 ;
      RECT  0.885000  0.645000  1.215000 1.030000 ;
      RECT  0.975000  1.030000  2.465000 1.215000 ;
      RECT  1.355000  2.630000  1.615000 2.905000 ;
      RECT  1.355000  2.905000  3.190000 3.075000 ;
      RECT  1.785000  0.085000  2.115000 0.860000 ;
      RECT  1.785000  2.460000  2.115000 2.735000 ;
      RECT  2.295000  0.580000  2.850000 0.860000 ;
      RECT  2.295000  1.215000  2.465000 2.905000 ;
      RECT  2.635000  0.860000  2.850000 2.735000 ;
      RECT  3.020000  2.035000  3.690000 2.375000 ;
      RECT  3.020000  2.375000  5.935000 2.545000 ;
      RECT  3.020000  2.545000  3.190000 2.905000 ;
      RECT  3.360000  2.715000  3.610000 3.245000 ;
      RECT  3.520000  0.295000  4.540000 0.465000 ;
      RECT  3.520000  0.465000  3.690000 2.035000 ;
      RECT  3.870000  0.635000  4.200000 2.035000 ;
      RECT  3.870000  2.035000  5.145000 2.205000 ;
      RECT  4.370000  0.465000  4.540000 1.335000 ;
      RECT  4.370000  1.335000  6.325000 1.505000 ;
      RECT  4.415000  2.715000  4.745000 3.245000 ;
      RECT  4.710000  0.085000  5.040000 1.165000 ;
      RECT  4.815000  1.675000  6.795000 1.845000 ;
      RECT  4.815000  1.845000  5.145000 2.035000 ;
      RECT  5.035000  2.715000  5.365000 2.905000 ;
      RECT  5.035000  2.905000  6.955000 3.075000 ;
      RECT  5.400000  2.015000  6.445000 2.205000 ;
      RECT  5.605000  2.545000  5.935000 2.735000 ;
      RECT  5.635000  0.265000  6.825000 0.435000 ;
      RECT  5.635000  0.435000  5.920000 0.965000 ;
      RECT  6.090000  0.645000  6.325000 1.335000 ;
      RECT  6.115000  2.205000  6.445000 2.735000 ;
      RECT  6.495000  0.435000  6.825000 0.855000 ;
      RECT  6.625000  1.845000  6.795000 2.365000 ;
      RECT  6.625000  2.365000  9.875000 2.535000 ;
      RECT  6.625000  2.705000  6.955000 2.905000 ;
      RECT  6.995000  0.255000  7.395000 0.640000 ;
      RECT  6.995000  0.640000  7.760000 0.970000 ;
      RECT  6.995000  0.970000  7.175000 1.940000 ;
      RECT  6.995000  1.940000  7.515000 2.195000 ;
      RECT  7.590000  1.565000  9.050000 1.735000 ;
      RECT  7.590000  1.735000  8.650000 1.770000 ;
      RECT  7.810000  2.705000  8.140000 3.245000 ;
      RECT  7.930000  0.085000  8.180000 0.970000 ;
      RECT  8.320000  1.770000  8.650000 2.195000 ;
      RECT  8.350000  0.640000  9.050000 0.970000 ;
      RECT  8.720000  0.970000  9.050000 1.565000 ;
      RECT  9.615000  0.660000  9.875000 2.365000 ;
      RECT  9.615000  2.535000  9.875000 2.775000 ;
      RECT 10.045000  0.660000 10.360000 1.380000 ;
      RECT 10.045000  1.380000 11.510000 1.550000 ;
      RECT 10.045000  1.550000 10.360000 2.775000 ;
      RECT 10.610000  1.720000 10.940000 1.795000 ;
      RECT 10.610000  1.795000 11.940000 1.975000 ;
      RECT 10.915000  2.145000 11.390000 3.245000 ;
      RECT 11.010000  0.085000 11.340000 1.210000 ;
      RECT 11.180000  1.550000 11.510000 1.625000 ;
      RECT 11.520000  0.590000 11.940000 1.210000 ;
      RECT 11.560000  1.975000 11.940000 2.375000 ;
      RECT 11.560000  2.375000 13.320000 2.545000 ;
      RECT 11.560000  2.545000 11.940000 2.755000 ;
      RECT 11.690000  1.210000 11.940000 1.795000 ;
      RECT 12.140000  0.085000 12.470000 0.880000 ;
      RECT 12.160000  2.715000 12.490000 3.245000 ;
      RECT 12.505000  1.405000 13.855000 1.585000 ;
      RECT 12.505000  1.585000 13.320000 1.655000 ;
      RECT 13.020000  2.715000 13.350000 3.245000 ;
      RECT 13.040000  0.085000 13.385000 1.140000 ;
      RECT 13.150000  1.655000 13.320000 2.375000 ;
      RECT 13.545000  1.755000 14.375000 1.925000 ;
      RECT 13.545000  1.925000 13.875000 2.485000 ;
      RECT 13.555000  0.325000 13.855000 1.055000 ;
      RECT 13.555000  1.055000 14.375000 1.225000 ;
      RECT 14.025000  1.225000 14.375000 1.755000 ;
      RECT 14.045000  0.085000 14.375000 0.885000 ;
      RECT 14.125000  2.105000 14.335000 3.245000 ;
      RECT 14.985000  0.085000 15.255000 1.090000 ;
      RECT 14.985000  1.815000 15.255000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
  END
END sky130_fd_sc_lp__sdfxbp_2
END LIBRARY
