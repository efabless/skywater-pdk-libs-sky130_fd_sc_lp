# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__or4bb_lp
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.405000 1.545000 5.865000 1.875000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.355000 1.815000 4.685000 2.150000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.400000 1.475000 1.795000 1.805000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.395000 1.110000 6.725000 1.780000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.265000 0.455000 0.595000 ;
        RECT 0.125000 0.595000 0.325000 2.325000 ;
        RECT 0.125000 2.325000 0.835000 3.065000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.505000  0.775000 1.595000 0.945000 ;
      RECT 0.505000  0.945000 0.675000 1.975000 ;
      RECT 0.505000  1.975000 1.220000 1.985000 ;
      RECT 0.505000  1.985000 2.365000 2.145000 ;
      RECT 0.855000  1.125000 1.945000 1.295000 ;
      RECT 0.855000  1.295000 1.130000 1.795000 ;
      RECT 0.915000  0.085000 1.245000 0.595000 ;
      RECT 1.035000  2.335000 1.365000 3.245000 ;
      RECT 1.050000  2.145000 2.365000 2.155000 ;
      RECT 1.425000  0.265000 2.035000 0.595000 ;
      RECT 1.425000  0.595000 1.595000 0.775000 ;
      RECT 1.565000  2.155000 2.365000 2.485000 ;
      RECT 1.565000  2.485000 1.895000 3.065000 ;
      RECT 1.775000  0.775000 3.200000 0.945000 ;
      RECT 1.775000  0.945000 1.945000 1.125000 ;
      RECT 2.035000  1.815000 2.365000 1.985000 ;
      RECT 2.360000  1.125000 2.690000 1.465000 ;
      RECT 2.360000  1.465000 2.715000 1.635000 ;
      RECT 2.505000  2.760000 2.835000 2.865000 ;
      RECT 2.505000  2.865000 5.155000 3.035000 ;
      RECT 2.545000  1.635000 2.715000 2.410000 ;
      RECT 2.545000  2.410000 4.175000 2.580000 ;
      RECT 2.870000  0.605000 3.200000 0.775000 ;
      RECT 2.870000  0.945000 3.200000 1.115000 ;
      RECT 2.870000  1.115000 4.340000 1.285000 ;
      RECT 3.495000  1.285000 3.825000 2.230000 ;
      RECT 3.660000  0.085000 3.990000 0.935000 ;
      RECT 4.005000  1.465000 5.035000 1.635000 ;
      RECT 4.005000  1.635000 4.175000 2.410000 ;
      RECT 4.170000  0.895000 4.780000 1.065000 ;
      RECT 4.170000  1.065000 4.340000 1.115000 ;
      RECT 4.355000  2.355000 4.685000 2.405000 ;
      RECT 4.355000  2.405000 6.725000 2.575000 ;
      RECT 4.355000  2.575000 4.685000 2.685000 ;
      RECT 4.450000  0.605000 4.780000 0.895000 ;
      RECT 4.865000  1.635000 5.035000 2.055000 ;
      RECT 4.865000  2.055000 6.215000 2.225000 ;
      RECT 5.320000  0.085000 5.650000 1.365000 ;
      RECT 5.830000  0.905000 6.215000 1.365000 ;
      RECT 5.845000  2.755000 6.175000 3.245000 ;
      RECT 5.965000  0.085000 6.295000 0.675000 ;
      RECT 6.045000  1.365000 6.215000 2.055000 ;
      RECT 6.395000  2.075000 7.085000 2.245000 ;
      RECT 6.395000  2.245000 6.725000 2.405000 ;
      RECT 6.395000  2.575000 6.725000 3.065000 ;
      RECT 6.755000  0.265000 7.085000 0.675000 ;
      RECT 6.915000  0.675000 7.085000 2.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_lp__or4bb_lp
END LIBRARY
