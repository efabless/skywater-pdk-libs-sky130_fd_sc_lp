# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__mux4_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.225000 1.580000 6.565000 1.910000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.475000 1.185000 4.680000 1.750000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.835000 1.485000 8.265000 2.860000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.765000 1.580000 7.045000 1.910000 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  0.477000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.795000 0.470000 8.985000 1.795000 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075000 1.185000 2.245000 2.120000 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.815000 1.645000 4.165000 1.815000 ;
        RECT 2.815000 1.815000 3.865000 1.985000 ;
        RECT 2.965000 0.360000 3.175000 0.860000 ;
        RECT 2.965000 0.860000 4.035000 1.030000 ;
        RECT 3.825000 0.360000 4.035000 0.860000 ;
        RECT 3.865000 1.030000 4.035000 1.210000 ;
        RECT 3.865000 1.210000 4.165000 1.645000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.600000 0.085000 ;
      RECT 0.000000  3.245000 9.600000 3.415000 ;
      RECT 0.155000  0.470000 0.365000 2.660000 ;
      RECT 0.605000  0.290000 2.375000 0.460000 ;
      RECT 0.605000  0.460000 0.795000 2.660000 ;
      RECT 1.035000  0.640000 1.245000 2.370000 ;
      RECT 1.035000  2.370000 4.215000 2.540000 ;
      RECT 1.035000  2.540000 1.245000 2.670000 ;
      RECT 1.425000  1.150000 1.895000 1.820000 ;
      RECT 1.565000  1.820000 1.895000 2.190000 ;
      RECT 1.725000  0.640000 2.025000 0.970000 ;
      RECT 1.725000  0.970000 1.895000 1.150000 ;
      RECT 2.205000  0.460000 2.375000 0.835000 ;
      RECT 2.205000  0.835000 2.785000 1.005000 ;
      RECT 2.325000  2.725000 2.655000 3.245000 ;
      RECT 2.555000  0.085000 2.745000 0.545000 ;
      RECT 2.615000  1.005000 2.785000 1.265000 ;
      RECT 2.615000  1.265000 3.640000 1.435000 ;
      RECT 3.185000  2.725000 3.515000 3.245000 ;
      RECT 3.395000  0.085000 3.605000 0.545000 ;
      RECT 4.045000  1.995000 5.075000 2.165000 ;
      RECT 4.045000  2.165000 4.215000 2.370000 ;
      RECT 4.255000  0.085000 4.465000 0.885000 ;
      RECT 4.395000  2.345000 4.725000 3.245000 ;
      RECT 4.905000  0.625000 5.345000 0.955000 ;
      RECT 4.905000  0.955000 5.075000 1.995000 ;
      RECT 4.905000  2.165000 5.075000 2.440000 ;
      RECT 4.905000  2.440000 5.600000 2.770000 ;
      RECT 5.255000  1.135000 5.695000 1.305000 ;
      RECT 5.255000  1.305000 5.425000 2.090000 ;
      RECT 5.255000  2.090000 7.620000 2.260000 ;
      RECT 5.525000  0.880000 7.525000 0.905000 ;
      RECT 5.525000  0.905000 6.645000 1.050000 ;
      RECT 5.525000  1.050000 5.695000 1.135000 ;
      RECT 5.605000  1.485000 6.045000 1.815000 ;
      RECT 5.875000  1.230000 8.615000 1.295000 ;
      RECT 5.875000  1.295000 7.655000 1.400000 ;
      RECT 5.875000  1.400000 6.045000 1.485000 ;
      RECT 5.965000  0.085000 6.295000 0.700000 ;
      RECT 6.270000  2.485000 6.600000 3.245000 ;
      RECT 6.475000  0.735000 7.525000 0.880000 ;
      RECT 7.230000  0.470000 7.525000 0.735000 ;
      RECT 7.410000  2.260000 7.620000 2.760000 ;
      RECT 7.485000  1.125000 8.615000 1.230000 ;
      RECT 7.485000  1.400000 7.655000 1.795000 ;
      RECT 8.070000  0.085000 8.400000 0.845000 ;
      RECT 8.445000  1.295000 8.615000 1.975000 ;
      RECT 8.445000  1.975000 9.495000 2.145000 ;
      RECT 8.490000  2.425000 8.700000 3.245000 ;
      RECT 8.920000  2.145000 9.130000 2.745000 ;
      RECT 9.165000  0.765000 9.495000 1.975000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  0.470000 0.325000 0.640000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  0.470000 7.525000 0.640000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
    LAYER met1 ;
      RECT 0.095000 0.440000 0.385000 0.485000 ;
      RECT 0.095000 0.485000 7.585000 0.625000 ;
      RECT 0.095000 0.625000 0.385000 0.670000 ;
      RECT 7.295000 0.440000 7.585000 0.485000 ;
      RECT 7.295000 0.625000 7.585000 0.670000 ;
  END
END sky130_fd_sc_lp__mux4_4
END LIBRARY
