# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__dlclkp_lp
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN GATE
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.605000 1.270000 2.150000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.389700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.755000 0.265000 7.110000 0.675000 ;
        RECT 6.845000 1.920000 7.110000 3.065000 ;
        RECT 6.940000 0.675000 7.110000 1.920000 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  0.689000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 5.020000 1.455000 5.635000 1.785000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.095000  0.265000 0.425000 0.715000 ;
      RECT 0.095000  0.715000 2.420000 0.885000 ;
      RECT 0.095000  0.885000 0.265000 2.330000 ;
      RECT 0.095000  2.330000 0.475000 3.065000 ;
      RECT 0.445000  1.065000 1.810000 1.395000 ;
      RECT 0.675000  2.330000 1.005000 3.245000 ;
      RECT 0.885000  0.085000 1.215000 0.535000 ;
      RECT 1.480000  1.395000 1.810000 1.450000 ;
      RECT 1.640000  1.450000 2.710000 1.780000 ;
      RECT 1.640000  1.780000 1.810000 2.515000 ;
      RECT 1.640000  2.515000 4.980000 2.685000 ;
      RECT 1.785000  0.265000 2.770000 0.535000 ;
      RECT 2.075000  2.075000 3.600000 2.335000 ;
      RECT 2.090000  0.885000 2.420000 1.095000 ;
      RECT 2.600000  0.535000 2.770000 0.815000 ;
      RECT 2.600000  0.815000 3.630000 1.145000 ;
      RECT 2.920000  1.325000 4.140000 1.495000 ;
      RECT 2.920000  1.495000 3.250000 1.715000 ;
      RECT 3.045000  0.085000 3.375000 0.635000 ;
      RECT 3.180000  2.865000 3.510000 3.245000 ;
      RECT 3.430000  1.675000 3.790000 1.935000 ;
      RECT 3.430000  1.935000 3.600000 2.075000 ;
      RECT 3.780000  2.155000 4.140000 2.335000 ;
      RECT 3.810000  0.265000 4.195000 0.505000 ;
      RECT 3.810000  0.505000 4.840000 0.675000 ;
      RECT 3.810000  0.675000 3.980000 1.325000 ;
      RECT 3.970000  1.495000 4.140000 2.155000 ;
      RECT 4.160000  0.895000 4.490000 1.145000 ;
      RECT 4.320000  1.145000 4.490000 2.315000 ;
      RECT 4.320000  2.315000 4.980000 2.515000 ;
      RECT 4.650000  2.685000 4.980000 3.065000 ;
      RECT 4.670000  0.675000 4.840000 1.965000 ;
      RECT 4.670000  1.965000 6.275000 2.135000 ;
      RECT 5.065000  0.085000 5.395000 1.275000 ;
      RECT 5.180000  2.315000 5.510000 3.245000 ;
      RECT 5.710000  2.315000 6.655000 2.485000 ;
      RECT 5.710000  2.485000 6.040000 3.065000 ;
      RECT 5.885000  0.905000 6.760000 1.075000 ;
      RECT 5.885000  1.075000 6.215000 1.365000 ;
      RECT 5.945000  1.545000 6.275000 1.965000 ;
      RECT 5.965000  0.085000 6.295000 0.675000 ;
      RECT 6.240000  2.665000 6.570000 3.245000 ;
      RECT 6.485000  1.075000 6.760000 1.575000 ;
      RECT 6.485000  1.575000 6.655000 2.315000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_lp__dlclkp_lp
END LIBRARY
