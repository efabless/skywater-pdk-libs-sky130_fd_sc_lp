# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__dfxbp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.995000 1.125000 2.255000 2.120000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.720000 0.255000 9.955000 1.140000 ;
        RECT 9.735000 1.140000 9.955000 3.075000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.640000 0.885000 8.970000 3.075000 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.840000 0.470000 1.795000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.560000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.560000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.560000 0.085000 ;
      RECT  0.000000  3.245000 10.560000 3.415000 ;
      RECT  0.095000  0.085000  0.425000 0.670000 ;
      RECT  0.095000  2.280000  0.405000 3.245000 ;
      RECT  0.575000  1.930000  1.040000 2.100000 ;
      RECT  0.575000  2.100000  0.855000 2.950000 ;
      RECT  0.595000  0.330000  1.040000 0.720000 ;
      RECT  0.790000  0.720000  1.040000 1.930000 ;
      RECT  1.140000  2.295000  1.475000 2.300000 ;
      RECT  1.140000  2.300000  2.170000 2.470000 ;
      RECT  1.140000  2.470000  1.410000 2.965000 ;
      RECT  1.215000  0.640000  1.475000 2.295000 ;
      RECT  1.580000  2.640000  1.830000 3.245000 ;
      RECT  1.645000  0.085000  1.975000 0.955000 ;
      RECT  2.000000  2.470000  2.170000 2.905000 ;
      RECT  2.000000  2.905000  3.475000 3.075000 ;
      RECT  2.180000  0.625000  2.595000 0.955000 ;
      RECT  2.350000  2.300000  2.595000 2.630000 ;
      RECT  2.425000  0.955000  2.595000 2.300000 ;
      RECT  2.765000  0.640000  3.015000 1.555000 ;
      RECT  2.765000  1.555000  4.285000 1.725000 ;
      RECT  2.765000  1.725000  2.945000 2.405000 ;
      RECT  2.765000  2.405000  3.125000 2.735000 ;
      RECT  3.125000  1.895000  3.475000 2.155000 ;
      RECT  3.305000  2.155000  3.475000 2.235000 ;
      RECT  3.305000  2.235000  5.145000 2.405000 ;
      RECT  3.305000  2.405000  3.475000 2.905000 ;
      RECT  3.475000  0.085000  4.355000 0.835000 ;
      RECT  3.485000  1.005000  4.785000 1.175000 ;
      RECT  3.485000  1.175000  3.815000 1.385000 ;
      RECT  3.945000  2.575000  4.275000 3.245000 ;
      RECT  4.025000  1.355000  4.285000 1.555000 ;
      RECT  4.455000  1.175000  4.785000 2.065000 ;
      RECT  4.525000  0.585000  4.785000 1.005000 ;
      RECT  4.955000  1.175000  5.145000 2.235000 ;
      RECT  5.075000  0.640000  5.565000 0.975000 ;
      RECT  5.315000  0.975000  5.565000 1.145000 ;
      RECT  5.315000  1.145000  6.795000 1.315000 ;
      RECT  5.315000  1.315000  5.565000 2.705000 ;
      RECT  5.970000  0.085000  6.490000 0.975000 ;
      RECT  5.995000  1.505000  6.325000 1.985000 ;
      RECT  5.995000  1.985000  7.170000 2.165000 ;
      RECT  6.270000  2.335000  6.730000 3.245000 ;
      RECT  6.535000  1.315000  6.795000 1.815000 ;
      RECT  6.660000  0.355000  7.135000 0.545000 ;
      RECT  6.660000  0.545000  9.540000 0.715000 ;
      RECT  6.660000  0.715000  7.135000 0.975000 ;
      RECT  6.900000  2.165000  7.170000 3.075000 ;
      RECT  6.965000  0.975000  7.135000 1.255000 ;
      RECT  6.965000  1.255000  7.435000 1.515000 ;
      RECT  6.965000  1.515000  7.170000 1.985000 ;
      RECT  7.545000  0.895000  8.470000 1.085000 ;
      RECT  7.545000  1.815000  7.815000 1.830000 ;
      RECT  7.545000  1.830000  7.875000 2.485000 ;
      RECT  7.605000  1.085000  8.470000 1.625000 ;
      RECT  7.605000  1.625000  7.815000 1.815000 ;
      RECT  8.045000  1.815000  8.470000 3.245000 ;
      RECT  8.095000  0.085000  8.425000 0.375000 ;
      RECT  9.150000  0.085000  9.480000 0.375000 ;
      RECT  9.150000  1.820000  9.480000 3.245000 ;
      RECT  9.370000  0.715000  9.540000 1.320000 ;
      RECT  9.370000  1.320000  9.555000 1.650000 ;
      RECT 10.125000  0.085000 10.420000 1.125000 ;
      RECT 10.125000  1.815000 10.415000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
  END
END sky130_fd_sc_lp__dfxbp_2
END LIBRARY
