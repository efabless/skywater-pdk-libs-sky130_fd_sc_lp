# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__sdfrbp_lp
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  19.20000 BY  3.330000 ;
  SYMMETRY R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.780000 0.265000 3.235000 0.435000 ;
        RECT 1.780000 0.435000 2.110000 0.535000 ;
        RECT 3.005000 0.435000 3.235000 0.670000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.598500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.755000 0.265000 19.085000 3.065000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.598500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.445000 0.265000 16.830000 1.075000 ;
        RECT 16.500000 1.765000 16.830000 3.065000 ;
        RECT 16.660000 1.075000 16.830000 1.765000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.633000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  3.935000 2.290000  4.225000 2.335000 ;
        RECT  3.935000 2.335000 14.305000 2.475000 ;
        RECT  3.935000 2.475000  4.225000 2.520000 ;
        RECT  6.815000 2.290000  7.105000 2.335000 ;
        RECT  6.815000 2.475000  7.105000 2.520000 ;
        RECT 14.015000 2.290000 14.305000 2.335000 ;
        RECT 14.015000 2.475000 14.305000 2.520000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.335000 1.550000 3.685000 1.965000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.477000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.475000 1.180000 0.805000 2.150000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 15.430000 1.295000 15.760000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 19.200000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 19.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 19.200000 0.085000 ;
      RECT  0.000000  3.245000 19.200000 3.415000 ;
      RECT  0.125000  0.265000  0.455000 0.715000 ;
      RECT  0.125000  0.715000  2.680000 0.885000 ;
      RECT  0.125000  0.885000  0.295000 2.435000 ;
      RECT  0.125000  2.435000  0.500000 3.065000 ;
      RECT  0.945000  0.085000  1.275000 0.535000 ;
      RECT  0.960000  2.495000  1.290000 3.245000 ;
      RECT  0.985000  1.065000  2.015000 1.235000 ;
      RECT  0.985000  1.235000  1.155000 2.145000 ;
      RECT  0.985000  2.145000  3.575000 2.315000 ;
      RECT  1.335000  1.415000  1.505000 1.795000 ;
      RECT  1.335000  1.795000  3.155000 1.965000 ;
      RECT  1.685000  1.235000  2.015000 1.615000 ;
      RECT  2.075000  2.315000  2.405000 3.065000 ;
      RECT  2.295000  0.615000  2.680000 0.715000 ;
      RECT  2.475000  1.065000  3.585000 1.235000 ;
      RECT  2.475000  1.235000  2.725000 1.615000 ;
      RECT  2.895000  2.495000  3.225000 3.245000 ;
      RECT  2.905000  1.415000  3.155000 1.795000 ;
      RECT  3.405000  2.315000  3.575000 2.700000 ;
      RECT  3.405000  2.700000  4.545000 2.975000 ;
      RECT  3.415000  0.725000  4.000000 0.895000 ;
      RECT  3.415000  0.895000  3.585000 1.065000 ;
      RECT  3.480000  0.085000  3.650000 0.555000 ;
      RECT  3.830000  0.265000  4.210000 0.715000 ;
      RECT  3.830000  0.715000  4.000000 0.725000 ;
      RECT  3.865000  1.625000  4.195000 2.520000 ;
      RECT  4.100000  1.075000  4.350000 1.445000 ;
      RECT  4.180000  0.885000  5.770000 1.055000 ;
      RECT  4.180000  1.055000  4.350000 1.075000 ;
      RECT  4.375000  2.025000  5.325000 2.195000 ;
      RECT  4.375000  2.195000  4.545000 2.700000 ;
      RECT  4.380000  0.265000  6.740000 0.435000 ;
      RECT  4.380000  0.435000  4.710000 0.715000 ;
      RECT  4.530000  1.235000  5.675000 1.405000 ;
      RECT  4.530000  1.405000  4.860000 1.535000 ;
      RECT  4.715000  2.385000  6.540000 2.555000 ;
      RECT  4.715000  2.555000  4.905000 2.895000 ;
      RECT  5.075000  1.585000  5.325000 2.025000 ;
      RECT  5.470000  0.715000  6.390000 0.885000 ;
      RECT  5.505000  1.405000  5.675000 1.545000 ;
      RECT  5.505000  1.545000  7.810000 1.715000 ;
      RECT  5.505000  1.715000  5.675000 2.385000 ;
      RECT  5.855000  1.885000  7.810000 2.055000 ;
      RECT  5.855000  2.055000  6.155000 2.215000 ;
      RECT  5.860000  2.735000  6.190000 3.245000 ;
      RECT  6.185000  1.065000  9.585000 1.165000 ;
      RECT  6.185000  1.165000  8.240000 1.235000 ;
      RECT  6.185000  1.235000  6.515000 1.375000 ;
      RECT  6.370000  2.555000  6.540000 2.700000 ;
      RECT  6.370000  2.700000  7.460000 2.870000 ;
      RECT  6.570000  0.435000  6.740000 0.715000 ;
      RECT  6.570000  0.715000  7.670000 0.885000 ;
      RECT  6.755000  2.225000  7.085000 2.520000 ;
      RECT  6.995000  0.085000  7.245000 0.535000 ;
      RECT  7.210000  2.870000  7.460000 3.065000 ;
      RECT  7.480000  1.415000  7.810000 1.545000 ;
      RECT  7.500000  0.265000  8.590000 0.435000 ;
      RECT  7.500000  0.435000  7.670000 0.715000 ;
      RECT  7.640000  2.055000  7.810000 2.895000 ;
      RECT  7.640000  2.895000  8.590000 3.065000 ;
      RECT  7.850000  0.615000  8.240000 0.995000 ;
      RECT  7.850000  0.995000  9.585000 1.065000 ;
      RECT  7.990000  1.235000  8.240000 2.715000 ;
      RECT  8.420000  0.435000  8.590000 0.645000 ;
      RECT  8.420000  0.645000 10.095000 0.815000 ;
      RECT  8.420000  1.345000  9.235000 1.675000 ;
      RECT  8.420000  1.675000  8.590000 2.895000 ;
      RECT  8.865000  0.085000  9.195000 0.465000 ;
      RECT  8.895000  1.855000  9.225000 3.245000 ;
      RECT  9.415000  1.165000  9.585000 2.895000 ;
      RECT  9.415000  2.895000 10.285000 3.065000 ;
      RECT  9.765000  0.265000 10.095000 0.645000 ;
      RECT  9.765000  0.815000 10.095000 1.435000 ;
      RECT  9.765000  1.435000 10.900000 1.765000 ;
      RECT  9.765000  1.765000  9.935000 2.715000 ;
      RECT 10.115000  1.945000 11.610000 2.115000 ;
      RECT 10.115000  2.115000 10.285000 2.895000 ;
      RECT 10.465000  2.295000 10.715000 2.895000 ;
      RECT 10.465000  2.895000 12.315000 3.065000 ;
      RECT 10.620000  0.575000 10.950000 1.085000 ;
      RECT 10.620000  1.085000 11.250000 1.255000 ;
      RECT 10.930000  2.425000 11.960000 2.595000 ;
      RECT 10.930000  2.595000 11.260000 2.715000 ;
      RECT 11.080000  1.255000 11.250000 1.915000 ;
      RECT 11.080000  1.915000 11.610000 1.945000 ;
      RECT 11.130000  0.575000 11.960000 0.905000 ;
      RECT 11.360000  2.115000 11.610000 2.245000 ;
      RECT 11.790000  0.905000 11.960000 1.745000 ;
      RECT 11.790000  1.745000 13.050000 1.915000 ;
      RECT 11.790000  1.915000 11.960000 2.425000 ;
      RECT 11.985000  2.795000 12.315000 2.895000 ;
      RECT 12.140000  1.050000 14.140000 1.060000 ;
      RECT 12.140000  1.060000 12.860000 1.220000 ;
      RECT 12.140000  1.220000 12.470000 1.565000 ;
      RECT 12.140000  2.185000 12.415000 2.445000 ;
      RECT 12.140000  2.445000 13.470000 2.615000 ;
      RECT 12.180000  0.085000 12.510000 0.870000 ;
      RECT 12.495000  2.795000 12.825000 3.245000 ;
      RECT 12.595000  2.095000 13.400000 2.265000 ;
      RECT 12.690000  0.265000 15.250000 0.435000 ;
      RECT 12.690000  0.435000 13.020000 0.595000 ;
      RECT 12.690000  0.890000 14.140000 1.050000 ;
      RECT 12.720000  1.400000 14.490000 1.570000 ;
      RECT 12.720000  1.570000 13.050000 1.745000 ;
      RECT 13.140000  2.615000 13.470000 3.030000 ;
      RECT 13.230000  1.750000 14.690000 1.920000 ;
      RECT 13.230000  1.920000 13.400000 2.095000 ;
      RECT 13.665000  2.100000 14.275000 2.520000 ;
      RECT 13.890000  0.685000 14.140000 0.890000 ;
      RECT 13.930000  2.700000 14.180000 3.245000 ;
      RECT 14.055000  1.240000 14.490000 1.400000 ;
      RECT 14.320000  0.890000 16.185000 1.060000 ;
      RECT 14.320000  1.060000 14.490000 1.240000 ;
      RECT 14.360000  2.700000 14.690000 3.030000 ;
      RECT 14.500000  0.435000 15.250000 0.710000 ;
      RECT 14.520000  1.920000 14.690000 2.700000 ;
      RECT 14.685000  1.240000 15.250000 1.570000 ;
      RECT 14.920000  1.570000 15.250000 3.065000 ;
      RECT 15.710000  0.085000 16.040000 0.710000 ;
      RECT 15.710000  1.960000 16.040000 3.245000 ;
      RECT 16.015000  1.060000 16.185000 1.255000 ;
      RECT 16.015000  1.255000 16.345000 1.585000 ;
      RECT 17.060000  0.665000 17.390000 1.305000 ;
      RECT 17.060000  1.305000 18.575000 1.635000 ;
      RECT 17.060000  1.635000 17.390000 2.495000 ;
      RECT 17.965000  0.085000 18.295000 1.125000 ;
      RECT 17.965000  1.815000 18.295000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  2.320000  4.165000 2.490000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  2.320000  7.045000 2.490000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  2.320000 14.245000 2.490000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.245000 15.685000 3.415000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.245000 16.165000 3.415000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.245000 16.645000 3.415000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.245000 17.125000 3.415000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.245000 17.605000 3.415000 ;
      RECT 17.915000 -0.085000 18.085000 0.085000 ;
      RECT 17.915000  3.245000 18.085000 3.415000 ;
      RECT 18.395000 -0.085000 18.565000 0.085000 ;
      RECT 18.395000  3.245000 18.565000 3.415000 ;
      RECT 18.875000 -0.085000 19.045000 0.085000 ;
      RECT 18.875000  3.245000 19.045000 3.415000 ;
  END
END sky130_fd_sc_lp__sdfrbp_lp
END LIBRARY
