# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__nand4bb_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015000 0.775000 1.305000 1.445000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.465000 0.775000 0.845000 1.445000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.855000 1.210000 4.645000 1.435000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.435000 1.425000 6.085000 1.750000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  2.125200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.210000 0.595000 2.435000 1.035000 ;
        RECT 2.210000 1.035000 3.685000 1.205000 ;
        RECT 2.325000 1.740000 5.265000 1.775000 ;
        RECT 2.325000 1.775000 4.235000 1.920000 ;
        RECT 2.325000 1.920000 2.515000 3.075000 ;
        RECT 3.185000 1.920000 3.375000 3.075000 ;
        RECT 3.420000 1.205000 3.685000 1.605000 ;
        RECT 3.420000 1.605000 5.265000 1.740000 ;
        RECT 4.045000 1.920000 4.235000 3.075000 ;
        RECT 4.905000 1.775000 5.265000 1.920000 ;
        RECT 4.905000 1.920000 5.475000 3.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.085000  0.275000 0.490000 0.605000 ;
      RECT 0.085000  0.605000 0.295000 1.625000 ;
      RECT 0.085000  1.625000 1.135000 1.795000 ;
      RECT 0.085000  1.795000 0.390000 2.240000 ;
      RECT 0.560000  1.965000 0.795000 3.245000 ;
      RECT 0.660000  0.085000 0.990000 0.555000 ;
      RECT 0.965000  1.795000 1.135000 2.345000 ;
      RECT 0.965000  2.345000 2.155000 2.515000 ;
      RECT 1.160000  0.275000 1.645000 0.605000 ;
      RECT 1.305000  1.845000 1.815000 2.175000 ;
      RECT 1.475000  0.605000 1.645000 1.325000 ;
      RECT 1.475000  1.325000 1.815000 1.845000 ;
      RECT 1.815000  0.255000 3.875000 0.425000 ;
      RECT 1.815000  0.425000 2.015000 1.095000 ;
      RECT 1.825000  2.685000 2.155000 3.245000 ;
      RECT 1.985000  1.375000 3.250000 1.570000 ;
      RECT 1.985000  1.570000 2.155000 2.345000 ;
      RECT 2.605000  0.425000 3.875000 0.465000 ;
      RECT 2.605000  0.465000 2.935000 0.825000 ;
      RECT 2.685000  2.105000 3.015000 3.245000 ;
      RECT 3.115000  0.635000 4.825000 0.865000 ;
      RECT 3.545000  2.090000 3.875000 3.245000 ;
      RECT 4.065000  0.255000 5.185000 0.465000 ;
      RECT 4.405000  1.945000 4.735000 3.245000 ;
      RECT 4.995000  0.465000 5.185000 1.065000 ;
      RECT 4.995000  1.065000 6.115000 1.235000 ;
      RECT 5.355000  0.085000 5.685000 0.895000 ;
      RECT 5.645000  1.920000 5.975000 3.245000 ;
      RECT 5.855000  0.255000 6.115000 1.065000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_lp__nand4bb_2
END LIBRARY
