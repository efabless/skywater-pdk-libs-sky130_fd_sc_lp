# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__a22o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.310000 1.200000 6.115000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.770000 1.345000 5.100000 1.615000 ;
        RECT 4.770000 1.615000 6.615000 1.785000 ;
        RECT 6.285000 1.210000 6.615000 1.615000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.400000 1.200000 4.020000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.970000 1.345000 3.230000 1.615000 ;
        RECT 2.970000 1.615000 4.560000 1.785000 ;
        RECT 4.230000 1.345000 4.560000 1.615000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 0.325000 0.425000 1.045000 ;
        RECT 0.100000 1.045000 2.460000 1.215000 ;
        RECT 0.100000 1.215000 0.345000 1.755000 ;
        RECT 0.100000 1.755000 2.050000 1.925000 ;
        RECT 0.960000 1.925000 1.150000 3.075000 ;
        RECT 1.410000 0.255000 1.590000 1.045000 ;
        RECT 1.820000 1.925000 2.050000 3.075000 ;
        RECT 2.270000 0.255000 2.460000 1.045000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.460000  2.095000 0.790000 3.245000 ;
      RECT 0.515000  1.385000 2.800000 1.585000 ;
      RECT 0.910000  0.085000 1.240000 0.875000 ;
      RECT 1.320000  2.095000 1.650000 3.245000 ;
      RECT 1.770000  0.085000 2.100000 0.865000 ;
      RECT 2.220000  1.815000 2.460000 3.245000 ;
      RECT 2.630000  0.085000 2.960000 0.650000 ;
      RECT 2.630000  0.820000 5.765000 1.030000 ;
      RECT 2.630000  1.030000 2.800000 1.385000 ;
      RECT 2.630000  1.585000 2.800000 1.955000 ;
      RECT 2.630000  1.955000 4.295000 2.135000 ;
      RECT 2.705000  2.305000 3.035000 2.905000 ;
      RECT 2.705000  2.905000 4.795000 3.075000 ;
      RECT 3.130000  0.255000 4.275000 0.650000 ;
      RECT 3.205000  2.135000 3.395000 2.735000 ;
      RECT 3.565000  2.305000 3.895000 2.905000 ;
      RECT 4.065000  2.135000 4.295000 2.735000 ;
      RECT 4.445000  0.085000 4.775000 0.650000 ;
      RECT 4.465000  1.955000 6.625000 2.125000 ;
      RECT 4.465000  2.125000 4.795000 2.905000 ;
      RECT 4.965000  2.295000 5.295000 3.245000 ;
      RECT 5.005000  0.255000 6.165000 0.530000 ;
      RECT 5.005000  0.530000 5.315000 0.650000 ;
      RECT 5.465000  2.125000 5.695000 3.075000 ;
      RECT 5.485000  0.700000 5.765000 0.820000 ;
      RECT 5.865000  2.295000 6.195000 3.245000 ;
      RECT 5.935000  0.530000 6.165000 1.030000 ;
      RECT 6.335000  0.085000 6.625000 1.030000 ;
      RECT 6.365000  2.125000 6.625000 3.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_lp__a22o_4
END LIBRARY
