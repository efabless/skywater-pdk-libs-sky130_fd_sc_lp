# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__srdlstp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.96000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.955000 0.455000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.594300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.505000 0.265000 12.835000 3.075000 ;
    END
  END Q
  PIN SET_B
    ANTENNAGATEAREA  0.409000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.980000 0.255000 5.765000 0.425000 ;
        RECT 1.980000 0.425000 2.310000 0.475000 ;
        RECT 5.435000 0.425000 5.765000 0.560000 ;
        RECT 5.435000 0.560000 5.635000 0.670000 ;
    END
  END SET_B
  PIN SLEEP_B
    ANTENNAGATEAREA  0.598000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.685000 1.480000 11.055000 2.150000 ;
    END
  END SLEEP_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 8.285000 1.480000 8.615000 2.150000 ;
    END
  END GATE
  PIN KAPWR
    ANTENNADIFFAREA  1.520900 ;
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 2.675000 12.890000 2.945000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.960000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.960000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.960000 0.085000 ;
      RECT  0.000000  3.245000 12.960000 3.415000 ;
      RECT  0.095000  0.085000  0.345000 0.785000 ;
      RECT  0.105000  1.980000  0.855000 2.150000 ;
      RECT  0.105000  2.150000  0.435000 2.660000 ;
      RECT  0.525000  0.325000  0.855000 0.785000 ;
      RECT  0.640000  2.320000  0.970000 3.245000 ;
      RECT  0.685000  0.785000  0.855000 1.480000 ;
      RECT  0.685000  1.480000  1.130000 1.810000 ;
      RECT  0.685000  1.810000  0.855000 1.980000 ;
      RECT  1.045000  0.630000  1.470000 1.310000 ;
      RECT  1.150000  1.980000  1.470000 2.505000 ;
      RECT  1.150000  2.505000  3.015000 2.675000 ;
      RECT  1.150000  2.675000  1.400000 2.860000 ;
      RECT  1.300000  1.310000  1.470000 1.980000 ;
      RECT  1.610000  2.845000  1.940000 3.245000 ;
      RECT  1.640000  0.085000  1.810000 0.645000 ;
      RECT  1.640000  0.645000  2.165000 0.815000 ;
      RECT  1.835000  0.815000  2.165000 1.310000 ;
      RECT  2.145000  1.480000  2.515000 2.335000 ;
      RECT  2.345000  0.850000  2.690000 0.985000 ;
      RECT  2.345000  0.985000  3.160000 1.255000 ;
      RECT  2.345000  1.255000  2.515000 1.480000 ;
      RECT  2.685000  1.425000  3.500000 1.595000 ;
      RECT  2.685000  1.595000  2.855000 2.265000 ;
      RECT  2.685000  2.265000  3.015000 2.505000 ;
      RECT  2.685000  2.675000  3.015000 3.075000 ;
      RECT  2.880000  0.595000  3.500000 0.815000 ;
      RECT  3.025000  1.765000  3.355000 2.095000 ;
      RECT  3.185000  2.095000  3.355000 2.905000 ;
      RECT  3.185000  2.905000  4.400000 3.075000 ;
      RECT  3.330000  0.815000  3.500000 1.425000 ;
      RECT  3.590000  2.075000  3.920000 2.735000 ;
      RECT  3.670000  0.595000  4.740000 0.895000 ;
      RECT  3.670000  0.895000  3.840000 2.075000 ;
      RECT  4.070000  1.125000  4.400000 1.455000 ;
      RECT  4.230000  1.455000  4.400000 2.315000 ;
      RECT  4.230000  2.315000  8.090000 2.485000 ;
      RECT  4.230000  2.485000  4.400000 2.905000 ;
      RECT  4.570000  0.895000  4.740000 1.285000 ;
      RECT  4.570000  1.285000  5.310000 1.455000 ;
      RECT  4.615000  2.655000  5.155000 3.075000 ;
      RECT  4.640000  1.625000  4.970000 1.975000 ;
      RECT  4.640000  1.975000  7.750000 2.145000 ;
      RECT  5.015000  0.595000  5.265000 0.840000 ;
      RECT  5.015000  0.840000  5.650000 1.010000 ;
      RECT  5.140000  1.455000  7.410000 1.515000 ;
      RECT  5.140000  1.515000  7.250000 1.625000 ;
      RECT  5.480000  1.010000  5.650000 1.115000 ;
      RECT  5.480000  1.115000  6.640000 1.285000 ;
      RECT  5.560000  1.625000  5.890000 1.805000 ;
      RECT  5.935000  0.085000  6.185000 0.945000 ;
      RECT  6.390000  0.615000  6.640000 1.115000 ;
      RECT  6.810000  2.655000  7.140000 2.985000 ;
      RECT  6.820000  0.085000  7.150000 1.015000 ;
      RECT  7.080000  1.185000  7.410000 1.455000 ;
      RECT  7.420000  1.685000  7.750000 1.975000 ;
      RECT  7.580000  0.800000  8.205000 0.970000 ;
      RECT  7.580000  0.970000  7.750000 1.685000 ;
      RECT  7.875000  0.340000  8.205000 0.800000 ;
      RECT  7.920000  1.140000  9.395000 1.310000 ;
      RECT  7.920000  1.310000  8.090000 2.315000 ;
      RECT  8.050000  2.745000  8.430000 3.075000 ;
      RECT  8.260000  2.320000 10.505000 2.490000 ;
      RECT  8.260000  2.490000  8.430000 2.745000 ;
      RECT  8.425000  0.850000  8.755000 1.140000 ;
      RECT  8.600000  2.660000  8.995000 2.990000 ;
      RECT  9.065000  1.310000  9.395000 2.150000 ;
      RECT  9.245000  2.660000  9.940000 2.990000 ;
      RECT  9.715000  0.085000 10.045000 1.310000 ;
      RECT 10.255000  0.635000 10.595000 1.095000 ;
      RECT 10.255000  1.095000 10.505000 2.320000 ;
      RECT 10.255000  2.490000 10.505000 2.860000 ;
      RECT 11.055000  0.085000 11.305000 1.095000 ;
      RECT 11.310000  1.475000 12.335000 1.645000 ;
      RECT 11.310000  1.645000 11.640000 2.495000 ;
      RECT 11.485000  0.635000 11.815000 1.315000 ;
      RECT 11.485000  1.315000 12.335000 1.475000 ;
      RECT 12.005000  1.815000 12.335000 3.245000 ;
      RECT 12.075000  0.085000 12.325000 1.145000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  2.735000  5.125000 2.905000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  2.735000  7.045000 2.905000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  2.735000  8.965000 2.905000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  2.735000  9.445000 2.905000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
  END
END sky130_fd_sc_lp__srdlstp_1
END LIBRARY
