# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__or2b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.000000 1.415000 2.775000 1.760000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.875000 0.470000 1.545000 ;
    END
  END B_N
  PIN X
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.080000 0.865000 1.445000 1.045000 ;
        RECT 1.080000 1.045000 1.410000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.095000  0.290000 0.420000 0.525000 ;
      RECT 0.095000  0.525000 2.860000 0.695000 ;
      RECT 0.160000  1.715000 0.820000 1.885000 ;
      RECT 0.160000  1.885000 0.490000 2.210000 ;
      RECT 0.590000  0.085000 0.935000 0.355000 ;
      RECT 0.650000  0.695000 0.820000 1.715000 ;
      RECT 0.685000  2.055000 0.910000 3.245000 ;
      RECT 1.580000  1.155000 1.830000 1.930000 ;
      RECT 1.580000  1.930000 3.060000 2.100000 ;
      RECT 1.580000  2.270000 1.840000 3.245000 ;
      RECT 1.615000  0.865000 2.520000 1.125000 ;
      RECT 1.615000  1.125000 1.830000 1.155000 ;
      RECT 1.625000  0.085000 1.955000 0.355000 ;
      RECT 2.690000  0.695000 2.860000 1.075000 ;
      RECT 2.690000  1.075000 3.635000 1.245000 ;
      RECT 2.730000  2.100000 3.060000 2.260000 ;
      RECT 2.945000  1.245000 3.635000 1.525000 ;
      RECT 3.030000  0.085000 3.360000 0.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__or2b_2
END LIBRARY
