# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__dlclkp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.960000 1.130000 1.335000 1.390000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 0.255000 6.590000 3.075000 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.435000 1.460000 3.845000 1.760000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.120000  0.255000 0.405000 0.665000 ;
      RECT 0.120000  0.665000 1.255000 0.835000 ;
      RECT 0.120000  0.835000 0.455000 1.095000 ;
      RECT 0.120000  1.095000 0.290000 1.910000 ;
      RECT 0.120000  1.910000 0.460000 2.630000 ;
      RECT 0.120000  2.630000 1.320000 2.800000 ;
      RECT 0.460000  1.345000 0.720000 1.560000 ;
      RECT 0.460000  1.560000 1.675000 1.730000 ;
      RECT 0.575000  0.085000 0.905000 0.495000 ;
      RECT 0.640000  2.970000 0.970000 3.245000 ;
      RECT 1.070000  1.730000 1.240000 2.280000 ;
      RECT 1.070000  2.280000 1.825000 2.450000 ;
      RECT 1.075000  0.265000 2.530000 0.435000 ;
      RECT 1.075000  0.435000 1.255000 0.665000 ;
      RECT 1.150000  2.800000 1.320000 2.905000 ;
      RECT 1.150000  2.905000 2.165000 3.075000 ;
      RECT 1.420000  1.900000 2.025000 1.930000 ;
      RECT 1.420000  1.930000 3.400000 1.985000 ;
      RECT 1.420000  1.985000 4.705000 2.110000 ;
      RECT 1.505000  0.605000 1.955000 0.845000 ;
      RECT 1.505000  0.845000 1.675000 1.560000 ;
      RECT 1.545000  2.450000 1.825000 2.735000 ;
      RECT 1.855000  1.015000 2.190000 1.265000 ;
      RECT 1.855000  1.265000 2.025000 1.900000 ;
      RECT 1.995000  2.345000 5.045000 2.515000 ;
      RECT 1.995000  2.515000 2.165000 2.905000 ;
      RECT 2.205000  1.475000 3.235000 1.760000 ;
      RECT 2.360000  0.435000 2.530000 0.935000 ;
      RECT 2.360000  0.935000 2.730000 1.265000 ;
      RECT 2.560000  2.685000 2.890000 3.245000 ;
      RECT 2.700000  0.085000 2.890000 0.765000 ;
      RECT 3.025000  0.875000 4.365000 1.065000 ;
      RECT 3.025000  1.065000 3.235000 1.475000 ;
      RECT 3.070000  0.485000 3.400000 0.525000 ;
      RECT 3.070000  0.525000 4.705000 0.695000 ;
      RECT 3.070000  2.110000 4.705000 2.175000 ;
      RECT 3.335000  2.515000 3.665000 3.075000 ;
      RECT 4.035000  1.065000 4.365000 1.815000 ;
      RECT 4.440000  0.085000 4.770000 0.345000 ;
      RECT 4.535000  0.695000 4.705000 1.985000 ;
      RECT 4.660000  2.685000 4.990000 3.245000 ;
      RECT 4.875000  1.345000 5.735000 1.535000 ;
      RECT 4.875000  1.535000 5.045000 2.345000 ;
      RECT 5.215000  1.705000 6.195000 1.875000 ;
      RECT 5.215000  1.875000 5.550000 2.495000 ;
      RECT 5.345000  0.710000 5.675000 1.005000 ;
      RECT 5.345000  1.005000 6.195000 1.175000 ;
      RECT 5.775000  2.045000 6.195000 3.245000 ;
      RECT 5.865000  0.085000 6.195000 0.835000 ;
      RECT 5.945000  1.175000 6.195000 1.705000 ;
      RECT 6.760000  0.085000 7.055000 1.095000 ;
      RECT 6.785000  1.815000 7.055000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_lp__dlclkp_2
END LIBRARY
