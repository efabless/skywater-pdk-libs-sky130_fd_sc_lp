# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__a2111oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.845000 1.210000 7.700000 1.435000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.945000 1.375000 9.975000 1.545000 ;
        RECT 7.945000 1.545000 8.485000 1.760000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.950000 1.425000 5.675000 1.760000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.050000 1.425000 3.740000 1.760000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.490000 1.210000 1.840000 1.435000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  2.587200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.140000 0.870000 2.505000 1.040000 ;
        RECT 0.140000 1.040000 0.320000 1.705000 ;
        RECT 0.140000 1.705000 1.645000 1.875000 ;
        RECT 0.595000 0.255000 0.785000 0.870000 ;
        RECT 0.595000 1.875000 0.785000 2.735000 ;
        RECT 1.455000 0.255000 1.645000 0.870000 ;
        RECT 1.455000 1.875000 1.645000 2.735000 ;
        RECT 2.305000 1.040000 2.505000 1.085000 ;
        RECT 2.305000 1.085000 5.185000 1.255000 ;
        RECT 2.315000 0.255000 2.505000 0.870000 ;
        RECT 3.175000 0.255000 3.425000 1.085000 ;
        RECT 4.095000 0.255000 4.335000 1.085000 ;
        RECT 4.945000 0.255000 5.195000 0.870000 ;
        RECT 4.945000 0.870000 7.605000 1.040000 ;
        RECT 4.945000 1.040000 5.185000 1.085000 ;
        RECT 6.460000 0.595000 6.705000 0.870000 ;
        RECT 7.310000 0.595000 7.605000 0.870000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.095000  0.085000  0.425000 0.700000 ;
      RECT 0.095000  2.045000  0.425000 2.905000 ;
      RECT 0.095000  2.905000  3.865000 3.075000 ;
      RECT 0.955000  0.085000  1.285000 0.700000 ;
      RECT 0.955000  2.045000  1.285000 2.905000 ;
      RECT 1.815000  0.085000  2.145000 0.700000 ;
      RECT 1.815000  1.930000  2.145000 2.905000 ;
      RECT 2.315000  1.930000  5.675000 2.100000 ;
      RECT 2.315000  2.100000  2.505000 2.735000 ;
      RECT 2.675000  0.085000  3.005000 0.915000 ;
      RECT 2.675000  2.270000  3.005000 2.905000 ;
      RECT 3.175000  2.100000  3.365000 2.735000 ;
      RECT 3.535000  2.270000  3.865000 2.905000 ;
      RECT 3.595000  0.085000  3.925000 0.915000 ;
      RECT 4.055000  2.270000  4.385000 2.905000 ;
      RECT 4.055000  2.905000  6.035000 3.075000 ;
      RECT 4.505000  0.085000  4.775000 0.915000 ;
      RECT 4.555000  2.100000  5.675000 2.120000 ;
      RECT 4.555000  2.120000  4.785000 2.735000 ;
      RECT 4.955000  2.305000  5.175000 2.905000 ;
      RECT 5.345000  2.120000  5.675000 2.735000 ;
      RECT 5.365000  0.085000  5.695000 0.690000 ;
      RECT 5.845000  1.605000  7.775000 1.775000 ;
      RECT 5.845000  1.775000  6.035000 2.905000 ;
      RECT 5.965000  0.255000  8.060000 0.425000 ;
      RECT 5.965000  0.425000  6.290000 0.700000 ;
      RECT 6.205000  1.945000  6.535000 3.245000 ;
      RECT 6.705000  1.775000  6.895000 3.075000 ;
      RECT 6.875000  0.425000  7.140000 0.700000 ;
      RECT 7.065000  1.945000  7.395000 3.245000 ;
      RECT 7.565000  1.775000  7.775000 1.930000 ;
      RECT 7.565000  1.930000  8.845000 2.100000 ;
      RECT 7.565000  2.100000  7.895000 3.075000 ;
      RECT 7.870000  0.425000  8.060000 1.035000 ;
      RECT 7.870000  1.035000  9.850000 1.205000 ;
      RECT 8.065000  2.270000  8.395000 3.245000 ;
      RECT 8.230000  0.085000  8.560000 0.865000 ;
      RECT 8.565000  2.100000  8.845000 3.075000 ;
      RECT 8.655000  1.715000  9.775000 1.885000 ;
      RECT 8.655000  1.885000  8.845000 1.930000 ;
      RECT 8.730000  0.255000  8.920000 1.035000 ;
      RECT 9.015000  2.055000  9.345000 3.245000 ;
      RECT 9.090000  0.085000  9.420000 0.865000 ;
      RECT 9.515000  1.885000  9.775000 3.075000 ;
      RECT 9.590000  0.255000  9.850000 1.035000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_lp__a2111oi_4
END LIBRARY
