# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__dfbbn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.88000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.180000 2.085000 1.510000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.010000 0.265000 14.340000 0.925000 ;
        RECT 14.010000 0.925000 14.445000 1.095000 ;
        RECT 14.010000 1.785000 14.445000 1.955000 ;
        RECT 14.010000 1.955000 14.340000 3.065000 ;
        RECT 14.275000 1.095000 14.445000 1.785000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.080000 0.265000 12.410000 1.005000 ;
        RECT 12.150000 1.695000 12.410000 2.990000 ;
        RECT 12.240000 1.005000 12.410000 1.695000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.165000 1.180000 11.560000 1.510000 ;
    END
  END RESET_B
  PIN SET_B
    ANTENNAPARTIALMETALSIDEAREA  3.115000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.795000 1.470000 9.575000 1.800000 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.910000 0.435000 2.150000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 14.880000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 14.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.880000 0.085000 ;
      RECT  0.000000  3.245000 14.880000 3.415000 ;
      RECT  0.110000  0.085000  0.360000 0.725000 ;
      RECT  0.140000  2.385000  0.470000 3.245000 ;
      RECT  0.540000  0.265000  0.870000 0.725000 ;
      RECT  0.650000  0.725000  0.870000 1.300000 ;
      RECT  0.650000  1.300000  1.005000 3.065000 ;
      RECT  1.090000  0.575000  1.420000 1.000000 ;
      RECT  1.210000  1.000000  1.380000 1.875000 ;
      RECT  1.210000  1.875000  2.560000 2.045000 ;
      RECT  1.210000  2.045000  1.540000 2.905000 ;
      RECT  1.600000  0.085000  1.930000 1.000000 ;
      RECT  1.720000  2.225000  2.050000 3.245000 ;
      RECT  2.290000  2.305000  2.910000 2.475000 ;
      RECT  2.290000  2.475000  2.620000 2.685000 ;
      RECT  2.295000  1.480000  2.560000 1.875000 ;
      RECT  2.445000  0.575000  2.775000 1.130000 ;
      RECT  2.445000  1.130000  2.910000 1.300000 ;
      RECT  2.740000  1.300000  2.910000 2.305000 ;
      RECT  3.035000  0.500000  3.260000 0.950000 ;
      RECT  3.090000  0.950000  3.260000 2.225000 ;
      RECT  3.090000  2.225000  3.990000 2.395000 ;
      RECT  3.090000  2.395000  3.420000 2.685000 ;
      RECT  3.440000  1.055000  4.885000 1.225000 ;
      RECT  3.440000  1.225000  3.640000 1.760000 ;
      RECT  3.820000  1.405000  4.720000 1.575000 ;
      RECT  3.820000  1.575000  3.990000 2.225000 ;
      RECT  4.170000  1.755000  4.370000 2.310000 ;
      RECT  4.170000  2.310000  6.055000 2.480000 ;
      RECT  4.205000  0.085000  4.535000 0.875000 ;
      RECT  4.550000  1.575000  4.720000 1.960000 ;
      RECT  4.550000  1.960000  5.705000 2.130000 ;
      RECT  4.630000  2.660000  4.960000 3.245000 ;
      RECT  4.715000  0.265000  6.680000 0.435000 ;
      RECT  4.715000  0.435000  4.885000 1.055000 ;
      RECT  4.900000  1.405000  5.165000 1.780000 ;
      RECT  5.065000  0.615000  6.330000 0.785000 ;
      RECT  5.065000  0.785000  5.395000 0.960000 ;
      RECT  5.140000  2.480000  5.470000 2.755000 ;
      RECT  5.375000  1.475000  5.705000 1.960000 ;
      RECT  5.575000  0.965000  5.905000 1.125000 ;
      RECT  5.575000  1.125000  6.055000 1.295000 ;
      RECT  5.885000  1.295000  6.055000 1.435000 ;
      RECT  5.885000  1.435000  7.155000 1.605000 ;
      RECT  5.885000  1.605000  6.055000 2.310000 ;
      RECT  6.160000  0.785000  6.330000 0.945000 ;
      RECT  6.235000  1.875000  6.565000 3.245000 ;
      RECT  6.510000  0.435000  6.680000 1.085000 ;
      RECT  6.510000  1.085000  7.775000 1.255000 ;
      RECT  6.825000  1.605000  7.155000 1.735000 ;
      RECT  6.860000  0.085000  7.110000 0.905000 ;
      RECT  7.335000  1.255000  7.775000 1.675000 ;
      RECT  7.335000  1.675000  7.505000 2.895000 ;
      RECT  7.335000  2.895000  8.615000 3.065000 ;
      RECT  7.685000  2.120000  8.125000 2.715000 ;
      RECT  7.955000  0.575000  8.285000 1.120000 ;
      RECT  7.955000  1.120000  9.955000 1.290000 ;
      RECT  7.955000  1.290000  8.125000 2.120000 ;
      RECT  8.345000  1.700000  8.615000 2.895000 ;
      RECT  8.885000  2.040000  9.215000 2.200000 ;
      RECT  8.885000  2.200000 11.965000 2.370000 ;
      RECT  9.035000  0.085000  9.365000 0.940000 ;
      RECT  9.355000  2.550000  9.605000 3.245000 ;
      RECT  9.545000  0.265000 10.905000 0.435000 ;
      RECT  9.545000  0.435000  9.875000 0.940000 ;
      RECT  9.785000  1.290000  9.955000 1.345000 ;
      RECT  9.785000  1.345000 10.125000 1.675000 ;
      RECT  9.785000  2.370000 10.115000 3.000000 ;
      RECT 10.135000  0.615000 10.475000 1.165000 ;
      RECT 10.305000  1.165000 10.475000 2.200000 ;
      RECT 10.575000  2.550000 10.905000 3.245000 ;
      RECT 10.655000  0.435000 10.905000 0.650000 ;
      RECT 10.655000  0.830000 11.470000 1.000000 ;
      RECT 10.655000  1.000000 10.985000 1.690000 ;
      RECT 10.815000  1.690000 11.460000 2.020000 ;
      RECT 11.220000  0.265000 11.470000 0.830000 ;
      RECT 11.640000  2.550000 11.970000 3.245000 ;
      RECT 11.650000  0.085000 11.900000 1.000000 ;
      RECT 11.795000  1.185000 12.060000 1.515000 ;
      RECT 11.795000  1.515000 11.965000 2.200000 ;
      RECT 12.590000  0.085000 12.840000 1.095000 ;
      RECT 12.590000  1.690000 12.840000 3.245000 ;
      RECT 13.070000  0.635000 13.400000 1.275000 ;
      RECT 13.070000  1.275000 14.095000 1.605000 ;
      RECT 13.070000  1.605000 13.400000 2.495000 ;
      RECT 13.580000  0.085000 13.830000 1.095000 ;
      RECT 13.580000  1.815000 13.830000 3.245000 ;
      RECT 14.520000  0.085000 14.770000 0.745000 ;
      RECT 14.520000  2.135000 14.770000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  1.580000  5.125000 1.750000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  1.580000  8.965000 1.750000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
    LAYER met1 ;
      RECT 4.895000 1.550000 5.185000 1.595000 ;
      RECT 4.895000 1.595000 9.025000 1.735000 ;
      RECT 4.895000 1.735000 5.185000 1.780000 ;
      RECT 8.735000 1.550000 9.025000 1.595000 ;
      RECT 8.735000 1.735000 9.025000 1.780000 ;
  END
END sky130_fd_sc_lp__dfbbn_2
END LIBRARY
