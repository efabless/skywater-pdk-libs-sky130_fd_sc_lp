/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/


`ifndef SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_14_TIMING_V
`define SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_14_TIMING_V

/**
 * sleep_pargate_plv: ????.
 *
 * Verilog simulation timing model.
 */

`timescale 1ns / 1ps
`default_nettype none

`celldefine
module sky130_fd_sc_lp__sleep_pargate_plv_14 (
    VIRTPWR,
    SLEEP
);

    // Module ports
    output VIRTPWR;
    input  SLEEP  ;

    // Module supplies
    supply1 VPWR;
    supply1 VPB ;
    supply0 VNB ;

    // Local signals
    wire vgnd;

    //       Name       Output   Other arguments
    pulldown pulldown0 (vgnd   );
    bufif0   bufif00   (VIRTPWR, VPWR, SLEEP    );

specify
(SLEEP => VIRTPWR) = (0:0:0,0:0:0,0:0:0,0:0:0,0:0:0,0:0:0);
endspecify
endmodule
`endcelldefine

`default_nettype wire
`endif  // SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_14_TIMING_V
