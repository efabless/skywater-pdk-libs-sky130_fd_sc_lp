# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__o2111a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.945000 1.415000 4.780000 1.760000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.370000 1.075000 5.335000 1.245000 ;
        RECT 3.370000 1.245000 3.775000 1.750000 ;
        RECT 5.165000 1.245000 5.335000 1.325000 ;
        RECT 5.165000 1.325000 5.495000 1.585000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.770000 1.425000 2.375000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225000 1.425000 1.600000 1.645000 ;
        RECT 1.430000 1.645000 1.600000 1.950000 ;
        RECT 1.430000 1.950000 2.735000 2.120000 ;
        RECT 2.555000 1.425000 2.985000 1.595000 ;
        RECT 2.555000 1.595000 2.735000 1.950000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.210000 0.390000 1.605000 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.865000 0.255000 6.090000 1.065000 ;
        RECT 5.865000 1.065000 7.595000 1.235000 ;
        RECT 6.015000 1.755000 7.595000 1.925000 ;
        RECT 6.015000 1.925000 6.205000 3.075000 ;
        RECT 6.760000 0.255000 6.950000 1.065000 ;
        RECT 6.875000 1.925000 7.065000 3.075000 ;
        RECT 7.235000 1.235000 7.595000 1.755000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.120000  1.815000 1.250000 1.985000 ;
      RECT 0.120000  1.985000 0.380000 3.075000 ;
      RECT 0.130000  0.255000 1.250000 0.425000 ;
      RECT 0.130000  0.425000 0.390000 1.040000 ;
      RECT 0.550000  2.155000 0.880000 3.245000 ;
      RECT 0.560000  0.595000 0.890000 1.815000 ;
      RECT 1.050000  1.985000 1.250000 2.290000 ;
      RECT 1.050000  2.290000 3.545000 2.460000 ;
      RECT 1.050000  2.460000 1.275000 3.075000 ;
      RECT 1.060000  0.425000 1.250000 1.085000 ;
      RECT 1.060000  1.085000 3.180000 1.255000 ;
      RECT 1.420000  0.285000 1.750000 0.725000 ;
      RECT 1.420000  0.725000 2.680000 0.915000 ;
      RECT 1.445000  2.630000 1.775000 3.245000 ;
      RECT 1.920000  0.255000 3.520000 0.425000 ;
      RECT 1.920000  0.425000 2.250000 0.555000 ;
      RECT 1.945000  2.460000 3.545000 2.470000 ;
      RECT 1.945000  2.470000 2.180000 3.075000 ;
      RECT 2.350000  2.640000 2.680000 3.245000 ;
      RECT 2.375000  0.680000 2.680000 0.725000 ;
      RECT 2.850000  0.595000 3.180000 1.085000 ;
      RECT 2.850000  2.470000 3.545000 3.075000 ;
      RECT 2.905000  1.930000 5.300000 2.100000 ;
      RECT 2.905000  2.100000 3.545000 2.290000 ;
      RECT 3.350000  0.425000 3.520000 0.725000 ;
      RECT 3.350000  0.725000 4.330000 0.735000 ;
      RECT 3.350000  0.735000 5.260000 0.905000 ;
      RECT 3.690000  0.085000 3.935000 0.545000 ;
      RECT 3.715000  2.280000 4.840000 2.450000 ;
      RECT 3.715000  2.450000 3.940000 3.075000 ;
      RECT 4.105000  0.255000 4.330000 0.725000 ;
      RECT 4.110000  2.620000 4.440000 3.245000 ;
      RECT 4.500000  0.085000 4.830000 0.565000 ;
      RECT 4.610000  2.450000 4.840000 3.075000 ;
      RECT 4.970000  1.755000 5.845000 1.925000 ;
      RECT 4.970000  1.925000 5.300000 1.930000 ;
      RECT 5.000000  0.255000 5.260000 0.735000 ;
      RECT 5.010000  2.100000 5.300000 3.075000 ;
      RECT 5.430000  0.085000 5.695000 0.930000 ;
      RECT 5.515000  2.105000 5.845000 3.245000 ;
      RECT 5.675000  1.405000 7.055000 1.585000 ;
      RECT 5.675000  1.585000 5.845000 1.755000 ;
      RECT 6.260000  0.085000 6.590000 0.895000 ;
      RECT 6.375000  2.095000 6.705000 3.245000 ;
      RECT 7.120000  0.085000 7.450000 0.895000 ;
      RECT 7.235000  2.095000 7.565000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_lp__o2111a_4
END LIBRARY
