# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__dlrtp_lp
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.080000 2.970000 1.410000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.619500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  9.645000 0.265000 10.440000 1.095000 ;
        RECT 10.110000 1.095000 10.440000 3.065000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.504000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.790000 1.345000 8.120000 1.780000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.835000 2.150000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.560000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.560000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.560000 0.085000 ;
      RECT 0.000000  3.245000 10.560000 3.415000 ;
      RECT 0.115000  0.085000  0.445000 0.725000 ;
      RECT 0.115000  2.330000  0.445000 3.245000 ;
      RECT 0.905000  0.265000  2.150000 0.435000 ;
      RECT 0.905000  0.435000  1.235000 0.725000 ;
      RECT 0.905000  2.330000  1.235000 3.010000 ;
      RECT 1.065000  0.725000  1.235000 2.330000 ;
      RECT 1.465000  0.615000  1.800000 3.065000 ;
      RECT 1.980000  0.435000  2.150000 0.895000 ;
      RECT 1.980000  0.895000  2.310000 1.590000 ;
      RECT 1.980000  1.590000  3.320000 1.760000 ;
      RECT 2.375000  0.085000  2.705000 0.715000 ;
      RECT 2.405000  1.940000  2.735000 3.245000 ;
      RECT 3.150000  0.895000  3.760000 1.225000 ;
      RECT 3.150000  1.225000  3.320000 1.590000 ;
      RECT 3.165000  0.345000  3.495000 0.545000 ;
      RECT 3.165000  0.545000  4.110000 0.715000 ;
      RECT 3.500000  1.405000  4.110000 1.575000 ;
      RECT 3.500000  1.575000  3.750000 2.735000 ;
      RECT 3.500000  2.735000  5.765000 3.065000 ;
      RECT 3.940000  0.715000  4.110000 1.405000 ;
      RECT 3.980000  1.755000  4.310000 2.385000 ;
      RECT 3.980000  2.385000  5.765000 2.555000 ;
      RECT 4.290000  0.265000  5.435000 0.435000 ;
      RECT 4.290000  0.435000  4.620000 0.945000 ;
      RECT 4.490000  1.345000  7.550000 1.515000 ;
      RECT 4.490000  1.515000  4.740000 2.205000 ;
      RECT 4.835000  0.615000  5.085000 1.345000 ;
      RECT 4.955000  1.695000  6.820000 1.865000 ;
      RECT 4.955000  1.865000  5.285000 2.155000 ;
      RECT 5.265000  0.435000  5.435000 0.995000 ;
      RECT 5.265000  0.995000  6.495000 1.165000 ;
      RECT 5.515000  2.045000  5.765000 2.385000 ;
      RECT 5.655000  0.085000  5.985000 0.815000 ;
      RECT 5.945000  2.045000  6.275000 3.245000 ;
      RECT 6.165000  0.485000  6.495000 0.995000 ;
      RECT 6.490000  1.865000  6.820000 2.375000 ;
      RECT 6.675000  0.265000  7.425000 0.645000 ;
      RECT 6.675000  0.645000  9.245000 0.815000 ;
      RECT 6.675000  0.815000  7.005000 0.935000 ;
      RECT 7.080000  1.815000  7.410000 2.325000 ;
      RECT 7.080000  2.325000  9.060000 2.495000 ;
      RECT 7.080000  2.495000  7.410000 3.065000 ;
      RECT 7.220000  0.995000  8.895000 1.165000 ;
      RECT 7.220000  1.165000  7.550000 1.345000 ;
      RECT 7.590000  2.675000  7.840000 3.245000 ;
      RECT 7.915000  0.085000  8.245000 0.465000 ;
      RECT 8.300000  1.815000  9.245000 1.985000 ;
      RECT 8.300000  1.985000  8.630000 2.145000 ;
      RECT 8.565000  1.165000  8.895000 1.625000 ;
      RECT 8.810000  2.165000  9.060000 2.325000 ;
      RECT 8.810000  2.495000  9.060000 3.065000 ;
      RECT 9.075000  0.815000  9.245000 1.185000 ;
      RECT 9.075000  1.185000  9.465000 1.515000 ;
      RECT 9.075000  1.515000  9.245000 1.815000 ;
      RECT 9.290000  2.165000  9.620000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
  END
END sky130_fd_sc_lp__dlrtp_lp
END LIBRARY
