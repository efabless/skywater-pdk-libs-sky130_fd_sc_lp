# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__sdfrbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.92000 BY  3.330000 ;
  SYMMETRY R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.475000 0.780000 1.805000 1.525000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.475000 0.355000 12.820000 2.285000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.395000 0.355000 13.765000 1.175000 ;
        RECT 13.400000 1.855000 13.765000 3.075000 ;
        RECT 13.585000 1.175000 13.765000 1.855000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  3.455000 1.920000  3.745000 1.965000 ;
        RECT  3.455000 1.965000 10.465000 2.105000 ;
        RECT  3.455000 2.105000  3.745000 2.150000 ;
        RECT  7.775000 1.920000  8.065000 1.965000 ;
        RECT  7.775000 2.105000  8.065000 2.150000 ;
        RECT 10.175000 1.920000 10.465000 1.965000 ;
        RECT 10.175000 2.105000 10.465000 2.150000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 1.155000 2.860000 2.215000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555000 1.535000 1.305000 1.695000 ;
        RECT 0.555000 1.695000 2.385000 1.865000 ;
        RECT 2.070000 1.395000 2.385000 1.695000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.410000 1.200000 4.645000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.920000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 13.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.920000 0.085000 ;
      RECT  0.000000  3.245000 13.920000 3.415000 ;
      RECT  0.155000  0.485000  0.365000 0.905000 ;
      RECT  0.155000  0.905000  1.235000 1.235000 ;
      RECT  0.155000  1.235000  0.325000 2.035000 ;
      RECT  0.155000  2.035000  2.375000 2.215000 ;
      RECT  0.585000  0.085000  0.795000 0.685000 ;
      RECT  0.590000  2.215000  0.920000 3.075000 ;
      RECT  1.045000  0.255000  3.105000 0.425000 ;
      RECT  1.045000  0.425000  1.305000 0.735000 ;
      RECT  1.090000  2.435000  1.350000 3.245000 ;
      RECT  1.810000  2.385000  3.210000 2.415000 ;
      RECT  1.810000  2.415000  3.275000 2.450000 ;
      RECT  1.810000  2.450000  6.035000 2.620000 ;
      RECT  1.810000  2.620000  2.140000 3.075000 ;
      RECT  1.985000  0.595000  2.315000 0.815000 ;
      RECT  1.985000  0.815000  3.210000 0.985000 ;
      RECT  2.775000  0.425000  3.105000 0.645000 ;
      RECT  2.775000  2.790000  3.105000 3.245000 ;
      RECT  3.040000  0.985000  3.210000 2.385000 ;
      RECT  3.275000  0.085000  3.605000 0.655000 ;
      RECT  3.275000  2.620000  3.605000 3.075000 ;
      RECT  3.380000  1.950000  3.750000 2.280000 ;
      RECT  4.235000  1.950000  4.995000 2.215000 ;
      RECT  4.255000  0.670000  4.425000 0.860000 ;
      RECT  4.255000  0.860000  4.995000 1.030000 ;
      RECT  4.665000  0.085000  4.995000 0.690000 ;
      RECT  4.665000  2.790000  4.995000 3.245000 ;
      RECT  4.825000  1.030000  4.995000 1.345000 ;
      RECT  4.825000  1.345000  5.150000 1.425000 ;
      RECT  4.825000  1.425000  5.230000 1.595000 ;
      RECT  4.825000  1.595000  5.150000 1.715000 ;
      RECT  4.825000  1.715000  4.995000 1.950000 ;
      RECT  5.165000  1.885000  6.175000 1.970000 ;
      RECT  5.165000  1.970000  5.480000 2.215000 ;
      RECT  5.185000  0.680000  5.485000 1.085000 ;
      RECT  5.185000  1.085000  5.535000 1.130000 ;
      RECT  5.185000  1.130000  6.175000 1.175000 ;
      RECT  5.290000  1.175000  6.175000 1.235000 ;
      RECT  5.320000  1.740000  6.175000 1.885000 ;
      RECT  5.345000  1.235000  6.175000 1.295000 ;
      RECT  5.400000  1.295000  6.175000 1.740000 ;
      RECT  5.655000  0.085000  5.835000 0.960000 ;
      RECT  5.775000  2.155000  6.515000 2.325000 ;
      RECT  5.775000  2.325000  6.035000 2.450000 ;
      RECT  5.775000  2.620000  6.035000 2.685000 ;
      RECT  6.005000  0.255000  7.780000 0.425000 ;
      RECT  6.005000  0.425000  6.175000 1.130000 ;
      RECT  6.205000  2.495000  7.990000 2.525000 ;
      RECT  6.205000  2.525000  6.905000 2.775000 ;
      RECT  6.345000  0.700000  6.515000 2.155000 ;
      RECT  6.725000  0.650000  6.945000 0.980000 ;
      RECT  6.725000  0.980000  6.895000 2.335000 ;
      RECT  6.725000  2.335000  7.990000 2.495000 ;
      RECT  7.065000  1.110000  8.915000 1.295000 ;
      RECT  7.065000  1.295000  7.245000 2.155000 ;
      RECT  7.075000  2.695000  7.405000 3.245000 ;
      RECT  7.105000  1.060000  8.915000 1.110000 ;
      RECT  7.425000  1.465000  8.575000 1.650000 ;
      RECT  7.425000  1.650000  7.605000 2.335000 ;
      RECT  7.585000  2.525000  7.990000 2.685000 ;
      RECT  7.610000  0.425000  7.780000 0.720000 ;
      RECT  7.610000  0.720000  9.255000 0.890000 ;
      RECT  7.775000  1.820000  8.080000 2.165000 ;
      RECT  7.950000  0.085000  8.280000 0.550000 ;
      RECT  8.250000  1.875000  8.480000 3.245000 ;
      RECT  8.660000  1.875000  8.915000 2.920000 ;
      RECT  8.745000  1.295000  8.915000 1.875000 ;
      RECT  9.085000  0.890000  9.255000 1.090000 ;
      RECT  9.085000  1.090000  9.350000 1.950000 ;
      RECT  9.085000  1.950000  9.720000 2.260000 ;
      RECT  9.190000  2.495000 10.060000 2.920000 ;
      RECT  9.425000  0.330000  9.830000 0.935000 ;
      RECT  9.540000  2.260000  9.720000 2.320000 ;
      RECT  9.550000  0.935000  9.830000 1.515000 ;
      RECT  9.550000  1.515000 10.680000 1.685000 ;
      RECT  9.550000  1.685000 10.060000 1.725000 ;
      RECT  9.890000  1.725000 10.060000 2.495000 ;
      RECT 10.000000  0.995000 10.805000 1.165000 ;
      RECT 10.000000  1.165000 10.340000 1.345000 ;
      RECT 10.135000  0.085000 10.465000 0.610000 ;
      RECT 10.230000  1.870000 10.795000 2.200000 ;
      RECT 10.350000  2.545000 10.610000 3.245000 ;
      RECT 10.510000  1.345000 11.190000 1.515000 ;
      RECT 10.635000  0.725000 11.590000 0.975000 ;
      RECT 10.635000  0.975000 10.805000 0.995000 ;
      RECT 10.790000  2.370000 11.135000 2.920000 ;
      RECT 10.965000  1.685000 11.590000 1.855000 ;
      RECT 10.965000  1.855000 11.135000 2.370000 ;
      RECT 10.975000  1.145000 11.190000 1.345000 ;
      RECT 11.025000  0.510000 11.355000 0.725000 ;
      RECT 11.305000  2.025000 11.635000 3.245000 ;
      RECT 11.360000  0.975000 11.590000 1.685000 ;
      RECT 11.545000  0.085000 11.875000 0.555000 ;
      RECT 11.805000  1.615000 12.305000 2.285000 ;
      RECT 11.970000  2.455000 13.230000 2.625000 ;
      RECT 11.970000  2.625000 12.300000 3.075000 ;
      RECT 12.045000  0.280000 12.305000 1.615000 ;
      RECT 12.900000  2.795000 13.230000 3.245000 ;
      RECT 12.990000  0.085000 13.225000 1.175000 ;
      RECT 13.040000  1.345000 13.415000 1.675000 ;
      RECT 13.040000  1.675000 13.230000 2.455000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  1.950000  3.685000 2.120000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  1.950000  8.005000 2.120000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  1.950000 10.405000 2.120000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
  END
END sky130_fd_sc_lp__sdfrbp_1
END LIBRARY
