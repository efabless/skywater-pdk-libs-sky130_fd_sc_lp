# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__o22a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.650000 1.075000 6.055000 1.185000 ;
        RECT 4.650000 1.185000 6.625000 1.245000 ;
        RECT 4.650000 1.245000 4.980000 1.515000 ;
        RECT 5.850000 1.245000 6.625000 1.770000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.190000 1.425000 5.680000 1.760000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.860000 1.195000 4.440000 1.245000 ;
        RECT 2.860000 1.245000 3.285000 1.525000 ;
        RECT 3.035000 1.075000 4.440000 1.195000 ;
        RECT 4.110000 1.245000 4.440000 1.515000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.455000 1.415000 3.900000 1.760000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 1.715000 1.225000 ;
        RECT 0.085000 1.225000 0.505000 1.755000 ;
        RECT 0.085000 1.755000 2.340000 1.925000 ;
        RECT 0.625000 0.255000 0.815000 1.055000 ;
        RECT 1.290000 1.925000 1.480000 3.075000 ;
        RECT 1.485000 0.255000 1.715000 1.055000 ;
        RECT 2.150000 1.925000 2.340000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.125000  0.085000 0.455000 0.885000 ;
      RECT 0.775000  1.405000 2.680000 1.575000 ;
      RECT 0.790000  2.095000 1.120000 3.245000 ;
      RECT 0.985000  0.085000 1.315000 0.885000 ;
      RECT 1.650000  2.105000 1.980000 3.245000 ;
      RECT 1.885000  0.085000 2.125000 1.105000 ;
      RECT 2.295000  0.255000 4.205000 0.515000 ;
      RECT 2.295000  0.515000 2.465000 1.405000 ;
      RECT 2.510000  1.575000 2.680000 1.930000 ;
      RECT 2.510000  1.930000 5.645000 2.100000 ;
      RECT 2.545000  2.270000 2.875000 3.245000 ;
      RECT 2.635000  0.685000 4.675000 0.735000 ;
      RECT 2.635000  0.735000 6.505000 0.905000 ;
      RECT 2.635000  0.905000 2.865000 1.015000 ;
      RECT 3.045000  2.270000 3.275000 2.905000 ;
      RECT 3.045000  2.905000 4.205000 3.075000 ;
      RECT 3.445000  2.100000 3.775000 2.735000 ;
      RECT 3.945000  2.270000 4.205000 2.905000 ;
      RECT 4.380000  2.270000 4.710000 3.245000 ;
      RECT 4.385000  0.255000 4.675000 0.685000 ;
      RECT 4.845000  0.085000 5.175000 0.565000 ;
      RECT 4.885000  2.270000 5.145000 2.905000 ;
      RECT 4.885000  2.905000 6.005000 3.075000 ;
      RECT 5.315000  2.100000 5.645000 2.735000 ;
      RECT 5.345000  0.255000 5.575000 0.735000 ;
      RECT 5.745000  0.085000 6.075000 0.565000 ;
      RECT 5.815000  1.940000 6.005000 2.905000 ;
      RECT 6.175000  1.940000 6.505000 3.245000 ;
      RECT 6.225000  0.905000 6.505000 1.015000 ;
      RECT 6.245000  0.255000 6.505000 0.735000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_lp__o22a_4
END LIBRARY
