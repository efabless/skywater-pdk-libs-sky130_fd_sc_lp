# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__dfsbp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.96000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.915000 1.365000 2.245000 1.605000 ;
        RECT 1.915000 1.605000 2.595000 2.515000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.145000 0.375000 12.390000 3.075000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.225000 0.255000 10.465000 3.075000 ;
    END
  END Q_N
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.315000 1.845000 5.505000 2.205000 ;
        RECT 5.315000 2.205000 6.605000 2.490000 ;
        RECT 6.435000 2.490000 6.605000 2.905000 ;
        RECT 6.435000 2.905000 7.620000 3.075000 ;
        RECT 7.430000 1.765000 8.345000 2.095000 ;
        RECT 7.430000 2.095000 7.620000 2.905000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.485000 0.540000 2.120000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.960000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.960000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.960000 0.085000 ;
      RECT  0.000000  3.245000 12.960000 3.415000 ;
      RECT  0.185000  0.085000  0.450000 1.270000 ;
      RECT  0.190000  2.290000  0.520000 3.245000 ;
      RECT  0.620000  1.015000  2.410000 1.195000 ;
      RECT  0.620000  1.195000  1.675000 1.305000 ;
      RECT  0.690000  2.290000  0.950000 2.630000 ;
      RECT  0.720000  1.305000  1.675000 1.485000 ;
      RECT  0.720000  1.485000  0.950000 2.290000 ;
      RECT  0.720000  2.630000  0.950000 2.775000 ;
      RECT  0.720000  2.775000  1.215000 3.075000 ;
      RECT  0.955000  0.255000  1.550000 0.845000 ;
      RECT  1.215000  1.805000  1.545000 2.305000 ;
      RECT  1.215000  2.305000  1.745000 2.475000 ;
      RECT  1.480000  2.475000  1.745000 2.975000 ;
      RECT  1.730000  0.085000  2.060000 0.845000 ;
      RECT  2.030000  2.685000  2.360000 3.245000 ;
      RECT  2.240000  0.255000  3.645000 0.425000 ;
      RECT  2.240000  0.425000  2.410000 1.015000 ;
      RECT  2.580000  0.670000  2.815000 1.265000 ;
      RECT  2.580000  1.265000  2.945000 1.435000 ;
      RECT  2.640000  2.695000  2.945000 3.025000 ;
      RECT  2.765000  1.435000  2.945000 2.695000 ;
      RECT  2.985000  0.670000  3.295000 1.000000 ;
      RECT  3.115000  1.000000  3.295000 2.365000 ;
      RECT  3.115000  2.365000  3.995000 2.535000 ;
      RECT  3.115000  2.535000  3.375000 3.045000 ;
      RECT  3.465000  0.425000  3.645000 1.125000 ;
      RECT  3.465000  1.125000  4.425000 1.295000 ;
      RECT  3.465000  1.295000  3.655000 2.185000 ;
      RECT  3.815000  0.085000  4.075000 0.955000 ;
      RECT  3.825000  1.815000  5.145000 1.985000 ;
      RECT  3.825000  1.985000  3.995000 2.365000 ;
      RECT  3.840000  2.835000  4.675000 3.245000 ;
      RECT  3.965000  1.465000  4.795000 1.645000 ;
      RECT  4.175000  2.185000  4.345000 2.495000 ;
      RECT  4.175000  2.495000  5.145000 2.665000 ;
      RECT  4.255000  0.515000  5.145000 0.720000 ;
      RECT  4.255000  0.720000  4.425000 1.125000 ;
      RECT  4.595000  0.890000  4.795000 1.465000 ;
      RECT  4.650000  1.985000  5.145000 2.325000 ;
      RECT  4.845000  2.665000  5.145000 2.720000 ;
      RECT  4.845000  2.720000  5.730000 3.075000 ;
      RECT  4.975000  0.720000  5.145000 1.165000 ;
      RECT  4.975000  1.165000  6.195000 1.335000 ;
      RECT  4.975000  1.505000  5.845000 1.675000 ;
      RECT  4.975000  1.675000  5.145000 1.815000 ;
      RECT  5.410000  0.085000  5.740000 0.995000 ;
      RECT  5.675000  1.675000  5.845000 1.705000 ;
      RECT  5.675000  1.705000  6.410000 2.035000 ;
      RECT  5.910000  0.265000  7.740000 0.465000 ;
      RECT  5.910000  0.465000  6.170000 0.995000 ;
      RECT  5.985000  2.660000  6.265000 3.245000 ;
      RECT  6.025000  1.335000  6.195000 1.355000 ;
      RECT  6.025000  1.355000  6.910000 1.525000 ;
      RECT  6.365000  0.635000  8.260000 0.805000 ;
      RECT  6.365000  0.805000  6.665000 1.170000 ;
      RECT  6.650000  1.525000  6.910000 2.025000 ;
      RECT  6.785000  2.405000  7.250000 2.735000 ;
      RECT  6.835000  0.975000  7.250000 1.175000 ;
      RECT  7.080000  1.175000  7.250000 1.405000 ;
      RECT  7.080000  1.405000  9.655000 1.585000 ;
      RECT  7.080000  1.585000  7.250000 2.405000 ;
      RECT  7.790000  2.275000  8.085000 3.245000 ;
      RECT  7.930000  0.500000  8.260000 0.635000 ;
      RECT  8.025000  0.985000  9.570000 1.065000 ;
      RECT  8.025000  1.065000 10.005000 1.235000 ;
      RECT  8.255000  2.275000  8.695000 2.605000 ;
      RECT  8.525000  1.585000  9.655000 1.645000 ;
      RECT  8.525000  1.645000  8.695000 2.275000 ;
      RECT  8.720000  0.085000  9.050000 0.815000 ;
      RECT  9.200000  1.815000 10.005000 1.985000 ;
      RECT  9.200000  1.985000  9.530000 2.210000 ;
      RECT  9.240000  0.700000  9.570000 0.985000 ;
      RECT  9.725000  2.155000 10.055000 3.245000 ;
      RECT  9.765000  0.085000 10.055000 0.895000 ;
      RECT  9.835000  1.235000 10.005000 1.815000 ;
      RECT 10.635000  0.085000 10.980000 1.095000 ;
      RECT 10.645000  1.815000 10.980000 3.245000 ;
      RECT 11.150000  0.700000 11.480000 1.345000 ;
      RECT 11.150000  1.345000 11.975000 1.675000 ;
      RECT 11.150000  1.675000 11.465000 2.485000 ;
      RECT 11.670000  0.085000 11.975000 1.175000 ;
      RECT 11.670000  1.845000 11.975000 3.245000 ;
      RECT 12.560000  0.085000 12.860000 1.255000 ;
      RECT 12.560000  1.815000 12.860000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
  END
END sky130_fd_sc_lp__dfsbp_2
END LIBRARY
