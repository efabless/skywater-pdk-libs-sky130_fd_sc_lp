# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__o221ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.405000 1.075000 8.590000 1.210000 ;
        RECT 6.405000 1.210000 9.990000 1.245000 ;
        RECT 6.405000 1.245000 6.655000 1.515000 ;
        RECT 8.385000 1.245000 9.990000 1.520000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.825000 1.425000 8.215000 1.750000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.810000 1.400000 3.820000 1.615000 ;
        RECT 2.810000 1.615000 6.145000 1.785000 ;
        RECT 5.815000 1.295000 6.145000 1.615000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.225000 1.195000 5.645000 1.445000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.425000 2.290000 1.750000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  2.654400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.595000 0.865000 1.085000 ;
        RECT 0.535000 1.085000 2.640000 1.255000 ;
        RECT 1.285000 1.920000 2.640000 1.955000 ;
        RECT 1.285000 1.955000 8.180000 2.090000 ;
        RECT 1.285000 2.090000 1.465000 3.075000 ;
        RECT 1.535000 0.595000 1.865000 1.085000 ;
        RECT 2.145000 2.090000 8.180000 2.120000 ;
        RECT 2.145000 2.120000 7.320000 2.125000 ;
        RECT 2.145000 2.125000 2.335000 3.075000 ;
        RECT 2.460000 1.255000 2.640000 1.920000 ;
        RECT 4.225000 2.125000 7.320000 2.135000 ;
        RECT 4.225000 2.135000 4.555000 2.735000 ;
        RECT 5.085000 2.135000 5.415000 2.735000 ;
        RECT 6.395000 1.950000 8.180000 1.955000 ;
        RECT 6.990000 2.135000 7.320000 2.735000 ;
        RECT 7.850000 2.120000 8.180000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.105000  0.255000  2.315000 0.425000 ;
      RECT 0.105000  0.425000  0.365000 1.185000 ;
      RECT 0.785000  1.920000  1.115000 3.245000 ;
      RECT 1.035000  0.425000  1.365000 0.895000 ;
      RECT 1.645000  2.260000  1.975000 3.245000 ;
      RECT 2.035000  0.425000  2.315000 0.655000 ;
      RECT 2.035000  0.655000  3.195000 0.915000 ;
      RECT 2.505000  0.255000  6.390000 0.445000 ;
      RECT 2.505000  0.445000  3.695000 0.485000 ;
      RECT 2.505000  2.295000  2.835000 3.245000 ;
      RECT 2.810000  0.915000  3.195000 1.005000 ;
      RECT 2.810000  1.005000  5.845000 1.025000 ;
      RECT 2.810000  1.025000  4.045000 1.230000 ;
      RECT 3.005000  2.295000  4.055000 2.465000 ;
      RECT 3.005000  2.465000  3.195000 3.075000 ;
      RECT 3.365000  0.485000  3.695000 0.835000 ;
      RECT 3.365000  2.635000  3.695000 3.245000 ;
      RECT 3.865000  0.615000  4.115000 0.775000 ;
      RECT 3.865000  0.775000  5.845000 1.005000 ;
      RECT 3.865000  2.465000  4.055000 2.905000 ;
      RECT 3.865000  2.905000  5.845000 3.075000 ;
      RECT 4.285000  0.445000  5.355000 0.605000 ;
      RECT 4.725000  2.315000  4.915000 2.905000 ;
      RECT 5.515000  0.665000  5.845000 0.775000 ;
      RECT 5.585000  2.305000  5.845000 2.905000 ;
      RECT 6.050000  2.305000  6.380000 3.245000 ;
      RECT 6.060000  0.445000  6.390000 0.735000 ;
      RECT 6.060000  0.735000  8.970000 0.870000 ;
      RECT 6.060000  0.870000  9.900000 0.905000 ;
      RECT 6.060000  0.905000  6.290000 0.945000 ;
      RECT 6.560000  0.085000  6.890000 0.565000 ;
      RECT 6.560000  2.305000  6.820000 2.905000 ;
      RECT 6.560000  2.905000  8.575000 3.075000 ;
      RECT 7.060000  0.255000  7.250000 0.735000 ;
      RECT 7.420000  0.085000  7.750000 0.565000 ;
      RECT 7.490000  2.290000  7.680000 2.905000 ;
      RECT 7.920000  0.255000  8.110000 0.735000 ;
      RECT 8.280000  0.085000  8.610000 0.565000 ;
      RECT 8.385000  1.690000  9.470000 1.860000 ;
      RECT 8.385000  1.860000  8.575000 2.905000 ;
      RECT 8.745000  2.030000  9.075000 3.245000 ;
      RECT 8.760000  0.905000  9.900000 1.040000 ;
      RECT 8.780000  0.255000  8.970000 0.735000 ;
      RECT 9.140000  0.085000  9.470000 0.700000 ;
      RECT 9.245000  1.860000  9.470000 3.075000 ;
      RECT 9.640000  0.255000  9.900000 0.870000 ;
      RECT 9.640000  1.815000  9.935000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_lp__o221ai_4
END LIBRARY
