# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__o32ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.425000 1.210000 10.455000 1.495000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.185000 1.210000 8.215000 1.495000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.335000 5.655000 1.760000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.065000 1.425000 3.755000 1.760000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.375000 1.855000 1.760000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  2.352000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 1.930000 6.005000 2.100000 ;
        RECT 0.540000 2.100000 0.870000 2.735000 ;
        RECT 0.570000 0.595000 0.800000 1.005000 ;
        RECT 0.570000 1.005000 6.005000 1.165000 ;
        RECT 0.570000 1.165000 3.410000 1.175000 ;
        RECT 1.400000 2.100000 1.765000 2.735000 ;
        RECT 1.470000 0.595000 1.660000 1.005000 ;
        RECT 2.330000 0.595000 2.520000 1.005000 ;
        RECT 3.190000 0.615000 3.380000 0.995000 ;
        RECT 3.190000 0.995000 6.005000 1.005000 ;
        RECT 4.570000 2.100000 4.820000 2.735000 ;
        RECT 5.415000 2.100000 5.680000 2.735000 ;
        RECT 5.835000 1.165000 6.005000 1.930000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.560000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.560000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.560000 0.085000 ;
      RECT 0.000000  3.245000 10.560000 3.415000 ;
      RECT 0.110000  0.255000  3.880000 0.425000 ;
      RECT 0.110000  0.425000  0.400000 1.095000 ;
      RECT 0.110000  1.940000  0.370000 2.905000 ;
      RECT 0.110000  2.905000  2.125000 3.075000 ;
      RECT 0.970000  0.425000  1.300000 0.835000 ;
      RECT 1.040000  2.270000  1.230000 2.905000 ;
      RECT 1.830000  0.425000  2.160000 0.835000 ;
      RECT 1.935000  2.270000  3.915000 2.450000 ;
      RECT 1.935000  2.450000  2.125000 2.905000 ;
      RECT 2.295000  2.620000  2.625000 3.245000 ;
      RECT 2.690000  0.425000  3.880000 0.445000 ;
      RECT 2.690000  0.445000  3.020000 0.835000 ;
      RECT 2.795000  2.450000  2.985000 3.075000 ;
      RECT 3.155000  2.620000  3.485000 3.245000 ;
      RECT 3.550000  0.445000  3.880000 0.655000 ;
      RECT 3.550000  0.655000  6.345000 0.825000 ;
      RECT 3.655000  2.450000  3.915000 3.075000 ;
      RECT 4.090000  0.085000  4.420000 0.485000 ;
      RECT 4.105000  2.270000  4.375000 2.905000 ;
      RECT 4.105000  2.905000  7.875000 3.075000 ;
      RECT 4.590000  0.255000  4.920000 0.655000 ;
      RECT 4.990000  2.270000  5.245000 2.905000 ;
      RECT 5.090000  0.085000  5.420000 0.485000 ;
      RECT 5.590000  0.255000  6.235000 0.645000 ;
      RECT 5.590000  0.645000  6.345000 0.655000 ;
      RECT 5.850000  2.270000  6.120000 2.905000 ;
      RECT 6.175000  0.825000  6.345000 0.870000 ;
      RECT 6.175000  0.870000 10.170000 1.040000 ;
      RECT 6.290000  1.665000  9.710000 1.835000 ;
      RECT 6.290000  1.835000  6.545000 2.735000 ;
      RECT 6.405000  0.085000  6.745000 0.475000 ;
      RECT 6.715000  2.005000  6.975000 2.905000 ;
      RECT 6.915000  0.255000  7.140000 0.870000 ;
      RECT 7.145000  1.835000  7.410000 2.735000 ;
      RECT 7.310000  0.085000  7.940000 0.700000 ;
      RECT 7.580000  2.005000  7.875000 2.905000 ;
      RECT 8.110000  0.255000  8.380000 0.870000 ;
      RECT 8.120000  2.005000  8.450000 3.245000 ;
      RECT 8.550000  0.085000  8.880000 0.700000 ;
      RECT 8.620000  1.835000  8.810000 3.075000 ;
      RECT 8.980000  2.005000  9.310000 3.245000 ;
      RECT 9.050000  0.255000  9.240000 0.870000 ;
      RECT 9.410000  0.085000  9.740000 0.700000 ;
      RECT 9.480000  1.835000  9.710000 3.075000 ;
      RECT 9.880000  1.815000 10.170000 3.245000 ;
      RECT 9.910000  0.255000 10.170000 0.870000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
  END
END sky130_fd_sc_lp__o32ai_4
END LIBRARY
