# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__ha_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.315000 1.570000 2.790000 1.760000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.885000 1.180000 2.145000 1.230000 ;
        RECT 1.885000 1.230000 3.270000 1.400000 ;
        RECT 1.885000 1.400000 2.145000 1.850000 ;
        RECT 2.960000 1.400000 3.270000 1.760000 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.325000 0.290000 4.715000 1.090000 ;
        RECT 4.395000 1.090000 4.715000 3.075000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.260000 0.365000 1.740000 ;
        RECT 0.095000 1.740000 0.505000 3.075000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.535000  0.085000 0.855000 1.060000 ;
      RECT 0.535000  1.230000 1.715000 1.400000 ;
      RECT 0.535000  1.400000 0.795000 1.560000 ;
      RECT 0.725000  1.815000 1.025000 3.245000 ;
      RECT 1.080000  0.355000 1.370000 1.230000 ;
      RECT 1.195000  1.600000 1.365000 2.675000 ;
      RECT 1.195000  2.675000 2.470000 2.885000 ;
      RECT 1.540000  0.355000 1.770000 0.840000 ;
      RECT 1.540000  0.840000 2.700000 1.010000 ;
      RECT 1.545000  1.400000 1.715000 2.175000 ;
      RECT 1.545000  2.175000 1.880000 2.505000 ;
      RECT 1.940000  0.085000 2.270000 0.670000 ;
      RECT 2.300000  1.930000 3.680000 2.100000 ;
      RECT 2.300000  2.100000 2.470000 2.675000 ;
      RECT 2.440000  0.355000 2.700000 0.840000 ;
      RECT 2.640000  2.270000 3.250000 3.245000 ;
      RECT 2.920000  0.755000 3.620000 1.060000 ;
      RECT 3.420000  2.100000 3.680000 2.505000 ;
      RECT 3.440000  1.060000 3.620000 1.260000 ;
      RECT 3.440000  1.260000 4.225000 1.590000 ;
      RECT 3.440000  1.590000 3.680000 1.930000 ;
      RECT 3.790000  0.085000 4.155000 1.090000 ;
      RECT 3.850000  1.815000 4.225000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_lp__ha_1
END LIBRARY
