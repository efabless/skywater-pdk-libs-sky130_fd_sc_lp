# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__mux2i_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.425000 1.715000 1.750000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.425000 1.335000 3.775000 1.760000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  1.575000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.435000 1.415000 7.045000 1.775000 ;
        RECT 4.435000 1.775000 9.025000 1.835000 ;
        RECT 6.875000 1.835000 9.025000 1.945000 ;
        RECT 8.855000 1.335000 9.170000 1.665000 ;
        RECT 8.855000 1.665000 9.025000 1.775000 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  2.961000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 0.325000 0.345000 1.075000 ;
        RECT 0.155000 1.075000 4.265000 1.165000 ;
        RECT 0.155000 1.165000 2.255000 1.245000 ;
        RECT 0.235000 1.930000 4.265000 2.100000 ;
        RECT 0.235000 2.100000 0.425000 2.940000 ;
        RECT 1.035000 0.635000 1.365000 0.965000 ;
        RECT 1.035000 0.965000 4.265000 1.075000 ;
        RECT 1.115000 2.100000 4.265000 2.110000 ;
        RECT 1.115000 2.110000 1.285000 2.600000 ;
        RECT 1.895000 1.245000 2.255000 1.470000 ;
        RECT 4.095000 1.165000 4.265000 1.930000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.600000 0.085000 ;
      RECT 0.000000  3.245000 9.600000 3.415000 ;
      RECT 0.525000  0.255000 1.795000 0.455000 ;
      RECT 0.525000  0.455000 0.855000 0.905000 ;
      RECT 0.665000  2.280000 0.875000 2.780000 ;
      RECT 0.665000  2.780000 1.735000 2.950000 ;
      RECT 1.525000  2.280000 6.615000 2.335000 ;
      RECT 1.525000  2.335000 4.615000 2.460000 ;
      RECT 1.525000  2.460000 1.735000 2.780000 ;
      RECT 1.535000  0.455000 1.795000 0.625000 ;
      RECT 1.535000  0.625000 4.615000 0.795000 ;
      RECT 2.385000  2.630000 7.565000 2.675000 ;
      RECT 2.385000  2.675000 4.965000 2.800000 ;
      RECT 2.385000  2.800000 3.455000 3.075000 ;
      RECT 2.405000  0.255000 4.965000 0.455000 ;
      RECT 4.445000  0.795000 4.615000 1.075000 ;
      RECT 4.445000  1.075000 8.335000 1.245000 ;
      RECT 4.445000  2.005000 6.615000 2.280000 ;
      RECT 4.795000  0.455000 4.965000 0.735000 ;
      RECT 4.795000  0.735000 6.685000 0.905000 ;
      RECT 4.795000  2.505000 7.565000 2.630000 ;
      RECT 4.940000  2.970000 5.270000 3.245000 ;
      RECT 5.135000  0.085000 5.325000 0.565000 ;
      RECT 5.495000  0.345000 5.825000 0.735000 ;
      RECT 5.915000  2.845000 6.245000 3.245000 ;
      RECT 5.995000  0.085000 6.185000 0.565000 ;
      RECT 6.355000  0.255000 6.685000 0.735000 ;
      RECT 6.795000  2.845000 7.125000 3.245000 ;
      RECT 6.855000  0.085000 7.115000 0.905000 ;
      RECT 6.880000  2.115000 8.575000 2.285000 ;
      RECT 6.880000  2.285000 7.565000 2.505000 ;
      RECT 7.225000  1.415000 8.675000 1.605000 ;
      RECT 7.285000  0.255000 7.475000 1.075000 ;
      RECT 7.295000  2.675000 7.565000 3.065000 ;
      RECT 7.645000  0.085000 7.975000 0.805000 ;
      RECT 7.735000  2.455000 8.065000 3.245000 ;
      RECT 8.145000  0.255000 8.335000 1.075000 ;
      RECT 8.235000  2.285000 8.575000 3.065000 ;
      RECT 8.505000  0.085000 8.835000 0.815000 ;
      RECT 8.505000  0.985000 9.510000 1.165000 ;
      RECT 8.505000  1.165000 8.675000 1.415000 ;
      RECT 8.745000  2.125000 9.025000 3.245000 ;
      RECT 9.005000  0.255000 9.205000 0.985000 ;
      RECT 9.195000  1.845000 9.510000 3.075000 ;
      RECT 9.340000  1.165000 9.510000 1.845000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
  END
END sky130_fd_sc_lp__mux2i_4
END LIBRARY
