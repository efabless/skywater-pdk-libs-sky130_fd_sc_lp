# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__bufbuf_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.48000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.355000 0.485000 1.750000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  4.704000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.625000 1.920000 11.935000 2.150000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.480000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.480000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.480000 0.085000 ;
      RECT  0.000000  3.245000 12.480000 3.415000 ;
      RECT  0.095000  0.255000  0.355000 1.015000 ;
      RECT  0.095000  1.015000  0.835000 1.185000 ;
      RECT  0.095000  1.920000  0.835000 2.090000 ;
      RECT  0.095000  2.090000  0.390000 3.075000 ;
      RECT  0.525000  0.085000  0.855000 0.845000 ;
      RECT  0.560000  2.260000  0.820000 3.245000 ;
      RECT  0.665000  1.185000  0.835000 1.405000 ;
      RECT  0.665000  1.405000  2.180000 1.590000 ;
      RECT  0.665000  1.590000  0.835000 1.920000 ;
      RECT  1.005000  1.760000  2.520000 1.930000 ;
      RECT  1.005000  1.930000  2.145000 1.945000 ;
      RECT  1.005000  1.945000  1.215000 3.075000 ;
      RECT  1.025000  0.255000  1.215000 1.065000 ;
      RECT  1.025000  1.065000  2.855000 1.235000 ;
      RECT  1.385000  0.085000  1.715000 0.895000 ;
      RECT  1.385000  2.115000  1.715000 3.245000 ;
      RECT  1.885000  0.255000  2.145000 1.065000 ;
      RECT  1.885000  1.945000  2.145000 3.075000 ;
      RECT  2.350000  1.235000  2.855000 1.385000 ;
      RECT  2.350000  1.385000  5.135000 1.575000 ;
      RECT  2.350000  1.575000  2.520000 1.760000 ;
      RECT  2.595000  0.085000  2.885000 0.895000 ;
      RECT  2.595000  2.100000  2.925000 3.245000 ;
      RECT  3.055000  0.255000  3.285000 1.045000 ;
      RECT  3.055000  1.045000  5.495000 1.215000 ;
      RECT  3.095000  1.745000  5.495000 1.925000 ;
      RECT  3.095000  1.925000  3.320000 3.075000 ;
      RECT  3.455000  0.085000  3.750000 0.875000 ;
      RECT  3.490000  2.095000  3.750000 3.245000 ;
      RECT  3.920000  0.255000  4.180000 1.045000 ;
      RECT  3.920000  1.925000  4.180000 3.075000 ;
      RECT  4.350000  0.085000  4.610000 0.875000 ;
      RECT  4.350000  2.095000  4.610000 3.245000 ;
      RECT  4.780000  0.255000  5.040000 1.045000 ;
      RECT  4.780000  1.925000  5.040000 3.075000 ;
      RECT  5.210000  0.085000  5.470000 0.875000 ;
      RECT  5.210000  2.095000  5.470000 3.245000 ;
      RECT  5.305000  1.215000  5.495000 1.745000 ;
      RECT  5.665000  0.255000  5.900000 3.075000 ;
      RECT  6.070000  0.085000  6.330000 1.075000 ;
      RECT  6.070000  1.315000  6.330000 1.755000 ;
      RECT  6.070000  1.925000  6.330000 3.245000 ;
      RECT  6.500000  0.255000  6.760000 3.075000 ;
      RECT  6.930000  0.085000  7.190000 1.075000 ;
      RECT  6.930000  1.315000  7.190000 1.755000 ;
      RECT  6.930000  1.925000  7.190000 3.245000 ;
      RECT  7.360000  0.255000  7.620000 3.075000 ;
      RECT  7.790000  0.085000  8.050000 1.075000 ;
      RECT  7.790000  1.315000  8.050000 1.755000 ;
      RECT  7.790000  1.925000  8.050000 3.245000 ;
      RECT  8.220000  0.255000  8.480000 3.075000 ;
      RECT  8.650000  0.085000  8.910000 1.075000 ;
      RECT  8.650000  1.315000  8.910000 1.755000 ;
      RECT  8.650000  1.925000  8.910000 3.245000 ;
      RECT  9.080000  0.255000  9.340000 3.075000 ;
      RECT  9.510000  0.085000  9.770000 1.075000 ;
      RECT  9.510000  1.315000  9.770000 1.755000 ;
      RECT  9.510000  1.925000  9.770000 3.245000 ;
      RECT  9.940000  0.255000 10.200000 3.075000 ;
      RECT 10.370000  0.085000 10.630000 1.075000 ;
      RECT 10.370000  1.315000 10.630000 1.755000 ;
      RECT 10.370000  1.925000 10.630000 3.245000 ;
      RECT 10.800000  0.255000 11.060000 3.075000 ;
      RECT 11.230000  0.085000 11.490000 1.075000 ;
      RECT 11.230000  1.315000 11.490000 1.755000 ;
      RECT 11.230000  1.925000 11.490000 3.245000 ;
      RECT 11.660000  0.255000 11.920000 3.075000 ;
      RECT 12.090000  0.085000 12.385000 1.075000 ;
      RECT 12.090000  1.925000 12.385000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.315000  1.580000  5.485000 1.750000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.685000  1.950000  5.855000 2.120000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.115000  1.580000  6.285000 1.750000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.545000  1.950000  6.715000 2.120000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  6.975000  1.580000  7.145000 1.750000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.405000  1.950000  7.575000 2.120000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  1.580000  8.005000 1.750000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.265000  1.950000  8.435000 2.120000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.695000  1.580000  8.865000 1.750000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.125000  1.950000  9.295000 2.120000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.555000  1.580000  9.725000 1.750000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT  9.985000  1.950000 10.155000 2.120000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.415000  1.580000 10.585000 1.750000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 10.845000  1.950000 11.015000 2.120000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.275000  1.580000 11.445000 1.750000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 11.705000  1.950000 11.875000 2.120000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
    LAYER met1 ;
      RECT 5.255000 1.550000 11.505000 1.780000 ;
  END
END sky130_fd_sc_lp__bufbuf_16
END LIBRARY
