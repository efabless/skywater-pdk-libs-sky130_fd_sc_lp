# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__fahcon_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.52000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.440000 1.345000 0.805000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.005000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.180000 5.050000 1.530000 ;
    END
  END B
  PIN CI
    ANTENNAGATEAREA  0.561000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.705000 1.180000 8.035000 1.515000 ;
    END
  END CI
  PIN COUT_N
    ANTENNADIFFAREA  1.035600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.875000 2.040000 6.205000 2.920000 ;
        RECT 6.035000 1.220000 6.475000 1.390000 ;
        RECT 6.035000 1.390000 6.205000 2.040000 ;
        RECT 6.305000 0.265000 6.635000 0.650000 ;
        RECT 6.305000 0.650000 6.475000 1.220000 ;
    END
  END COUT_N
  PIN SUM
    ANTENNADIFFAREA  0.579600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.155000 0.265000 11.420000 3.065000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.520000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.520000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.520000 0.085000 ;
      RECT  0.000000  3.245000 11.520000 3.415000 ;
      RECT  0.090000  0.375000  0.490000 0.995000 ;
      RECT  0.090000  0.995000  1.190000 1.165000 ;
      RECT  0.090000  1.165000  0.260000 1.960000 ;
      RECT  0.090000  1.960000  0.475000 3.065000 ;
      RECT  0.655000  1.960000  0.985000 3.245000 ;
      RECT  0.670000  0.085000  0.840000 0.815000 ;
      RECT  0.985000  1.345000  1.190000 1.675000 ;
      RECT  1.020000  0.265000  2.705000 0.435000 ;
      RECT  1.020000  0.435000  1.190000 0.995000 ;
      RECT  1.020000  1.165000  1.190000 1.345000 ;
      RECT  1.210000  1.855000  1.540000 2.895000 ;
      RECT  1.210000  2.895000  3.805000 3.065000 ;
      RECT  1.370000  0.615000  1.710000 1.235000 ;
      RECT  1.370000  1.235000  1.540000 1.855000 ;
      RECT  1.720000  1.415000  2.275000 1.585000 ;
      RECT  1.720000  1.585000  1.890000 2.545000 ;
      RECT  1.720000  2.545000  3.260000 2.715000 ;
      RECT  1.890000  0.615000  2.275000 1.415000 ;
      RECT  2.070000  1.775000  2.240000 2.195000 ;
      RECT  2.070000  2.195000  3.260000 2.365000 ;
      RECT  2.420000  1.765000  2.750000 2.015000 ;
      RECT  2.455000  0.435000  2.705000 1.765000 ;
      RECT  2.885000  0.265000  4.665000 0.435000 ;
      RECT  2.885000  0.435000  3.215000 0.525000 ;
      RECT  2.930000  0.705000  3.260000 2.195000 ;
      RECT  3.475000  0.615000  3.910000 1.295000 ;
      RECT  3.475000  1.295000  3.805000 2.895000 ;
      RECT  4.055000  1.775000  4.385000 3.065000 ;
      RECT  4.095000  0.435000  4.665000 1.000000 ;
      RECT  4.095000  1.000000  4.265000 1.775000 ;
      RECT  4.565000  1.775000  4.895000 3.245000 ;
      RECT  4.845000  0.085000  5.095000 1.000000 ;
      RECT  5.145000  1.880000  5.475000 2.920000 ;
      RECT  5.305000  0.460000  6.125000 0.630000 ;
      RECT  5.305000  0.630000  5.475000 1.880000 ;
      RECT  5.655000  0.810000  6.115000 1.040000 ;
      RECT  5.655000  1.040000  5.855000 1.740000 ;
      RECT  5.795000  0.265000  6.125000 0.460000 ;
      RECT  6.385000  1.570000  6.650000 2.150000 ;
      RECT  6.655000  0.830000  7.045000 1.330000 ;
      RECT  6.860000  1.510000  7.475000 1.680000 ;
      RECT  6.860000  1.680000  7.110000 2.920000 ;
      RECT  7.225000  0.265000  7.475000 1.510000 ;
      RECT  7.320000  1.860000  7.650000 3.245000 ;
      RECT  7.785000  0.085000  8.035000 1.000000 ;
      RECT  7.830000  1.815000  8.385000 2.545000 ;
      RECT  7.830000  2.545000 10.025000 2.715000 ;
      RECT  7.830000  2.715000  8.160000 3.065000 ;
      RECT  8.215000  0.265000  8.550000 1.045000 ;
      RECT  8.215000  1.045000  8.385000 1.815000 ;
      RECT  8.520000  2.895000 10.455000 3.065000 ;
      RECT  8.565000  1.225000  8.745000 1.725000 ;
      RECT  8.565000  1.725000  8.965000 1.895000 ;
      RECT  8.765000  0.265000 10.375000 0.435000 ;
      RECT  8.765000  0.435000  9.095000 1.045000 ;
      RECT  8.765000  1.895000  8.965000 2.150000 ;
      RECT  8.925000  1.045000  9.095000 1.220000 ;
      RECT  8.925000  1.220000  9.315000 1.390000 ;
      RECT  9.145000  1.390000  9.315000 2.365000 ;
      RECT  9.275000  0.810000  9.675000 1.040000 ;
      RECT  9.495000  1.040000  9.675000 1.855000 ;
      RECT  9.495000  2.035000 10.025000 2.545000 ;
      RECT  9.855000  0.615000 10.025000 1.075000 ;
      RECT  9.855000  1.075000 10.580000 1.245000 ;
      RECT  9.855000  1.425000 10.230000 1.755000 ;
      RECT  9.855000  1.755000 10.025000 2.035000 ;
      RECT 10.205000  0.435000 10.375000 0.725000 ;
      RECT 10.205000  0.725000 10.975000 0.895000 ;
      RECT 10.205000  1.935000 10.580000 2.105000 ;
      RECT 10.205000  2.105000 10.455000 2.895000 ;
      RECT 10.410000  1.245000 10.580000 1.935000 ;
      RECT 10.610000  0.085000 10.860000 0.545000 ;
      RECT 10.660000  2.285000 10.910000 3.245000 ;
      RECT 10.760000  0.895000 10.975000 1.515000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  0.840000  2.245000 1.010000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  1.950000  3.205000 2.120000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  0.840000  6.085000 1.010000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  1.950000  6.565000 2.120000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  0.840000  7.045000 1.010000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  1.950000  8.965000 2.120000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  0.840000  9.445000 1.010000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
    LAYER met1 ;
      RECT 2.015000 0.810000 2.305000 0.855000 ;
      RECT 2.015000 0.855000 9.505000 0.995000 ;
      RECT 2.015000 0.995000 2.305000 1.040000 ;
      RECT 2.975000 1.920000 3.265000 1.965000 ;
      RECT 2.975000 1.965000 9.025000 2.105000 ;
      RECT 2.975000 2.105000 3.265000 2.150000 ;
      RECT 5.855000 0.810000 6.145000 0.855000 ;
      RECT 5.855000 0.995000 6.145000 1.040000 ;
      RECT 6.335000 1.920000 6.625000 1.965000 ;
      RECT 6.335000 2.105000 6.625000 2.150000 ;
      RECT 6.815000 0.810000 7.105000 0.855000 ;
      RECT 6.815000 0.995000 7.105000 1.040000 ;
      RECT 8.735000 1.920000 9.025000 1.965000 ;
      RECT 8.735000 2.105000 9.025000 2.150000 ;
      RECT 9.215000 0.810000 9.505000 0.855000 ;
      RECT 9.215000 0.995000 9.505000 1.040000 ;
  END
END sky130_fd_sc_lp__fahcon_1
END LIBRARY
