# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__a22oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625000 1.345000 0.885000 1.950000 ;
        RECT 0.625000 1.950000 2.375000 2.120000 ;
        RECT 2.125000 1.345000 2.375000 1.950000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055000 1.345000 1.915000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905000 1.345000 3.155000 1.925000 ;
        RECT 2.905000 1.925000 4.165000 2.095000 ;
        RECT 3.985000 1.345000 4.555000 1.750000 ;
        RECT 3.985000 1.750000 4.165000 1.925000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365000 1.345000 3.815000 1.750000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.604400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.440000 0.255000 0.690000 0.995000 ;
        RECT 0.440000 0.995000 2.740000 1.005000 ;
        RECT 0.440000 1.005000 4.680000 1.165000 ;
        RECT 2.410000 0.255000 2.740000 0.995000 ;
        RECT 2.550000 1.165000 4.680000 1.175000 ;
        RECT 2.550000 1.175000 2.735000 2.265000 ;
        RECT 2.550000 2.265000 4.240000 2.435000 ;
        RECT 3.920000 2.435000 4.240000 2.595000 ;
        RECT 4.400000 0.255000 4.680000 1.005000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.205000  1.855000 0.455000 2.290000 ;
      RECT 0.205000  2.290000 2.380000 2.460000 ;
      RECT 0.205000  2.460000 0.535000 3.075000 ;
      RECT 0.750000  2.630000 1.080000 3.245000 ;
      RECT 0.870000  0.265000 1.200000 0.655000 ;
      RECT 0.870000  0.655000 2.220000 0.825000 ;
      RECT 1.280000  2.460000 1.540000 3.075000 ;
      RECT 1.380000  0.085000 1.710000 0.485000 ;
      RECT 1.710000  2.630000 2.040000 2.945000 ;
      RECT 1.710000  2.945000 2.410000 3.245000 ;
      RECT 1.890000  0.265000 2.220000 0.655000 ;
      RECT 2.210000  2.460000 2.380000 2.605000 ;
      RECT 2.210000  2.605000 3.725000 2.765000 ;
      RECT 2.210000  2.765000 4.680000 2.775000 ;
      RECT 2.590000  2.775000 4.680000 3.075000 ;
      RECT 2.980000  0.255000 3.320000 0.665000 ;
      RECT 2.980000  0.665000 4.230000 0.835000 ;
      RECT 3.490000  0.085000 3.820000 0.495000 ;
      RECT 3.990000  0.505000 4.230000 0.665000 ;
      RECT 4.410000  1.990000 4.680000 2.765000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_lp__a22oi_2
END LIBRARY
