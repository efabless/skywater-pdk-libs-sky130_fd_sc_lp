# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__o32a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.500000 1.210000 1.830000 1.525000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.425000 1.330000 1.695000 ;
        RECT 0.085000 1.695000 2.180000 1.865000 ;
        RECT 2.010000 1.270000 2.375000 1.535000 ;
        RECT 2.010000 1.535000 2.180000 1.695000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 1.210000 3.690000 1.535000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.210000 4.775000 1.525000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.860000 1.355000 4.195000 1.695000 ;
        RECT 3.860000 1.695000 5.625000 1.865000 ;
        RECT 4.945000 1.425000 5.625000 1.695000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.485000 0.255000 6.665000 1.055000 ;
        RECT 6.485000 1.055000 8.075000 1.225000 ;
        RECT 6.485000 1.755000 8.075000 1.925000 ;
        RECT 6.485000 1.925000 6.675000 3.075000 ;
        RECT 7.345000 0.255000 7.525000 1.055000 ;
        RECT 7.345000 1.925000 7.535000 3.075000 ;
        RECT 7.810000 1.225000 8.075000 1.755000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.180000  0.305000 0.440000 1.085000 ;
      RECT 0.180000  1.085000 1.330000 1.255000 ;
      RECT 0.520000  2.035000 2.540000 2.205000 ;
      RECT 0.520000  2.205000 0.780000 3.065000 ;
      RECT 0.610000  0.085000 1.235000 0.700000 ;
      RECT 0.610000  0.700000 0.940000 0.915000 ;
      RECT 0.950000  2.375000 2.180000 2.545000 ;
      RECT 0.950000  2.545000 1.210000 3.075000 ;
      RECT 1.160000  0.870000 3.855000 1.040000 ;
      RECT 1.160000  1.040000 1.330000 1.085000 ;
      RECT 1.380000  2.715000 1.710000 3.245000 ;
      RECT 1.405000  0.255000 1.640000 0.870000 ;
      RECT 1.810000  0.085000 2.140000 0.700000 ;
      RECT 1.880000  2.545000 2.180000 3.075000 ;
      RECT 2.310000  0.305000 2.560000 0.870000 ;
      RECT 2.350000  1.705000 3.470000 1.875000 ;
      RECT 2.350000  1.875000 2.540000 2.035000 ;
      RECT 2.350000  2.205000 2.540000 3.075000 ;
      RECT 2.710000  2.045000 3.040000 2.905000 ;
      RECT 2.710000  2.905000 3.920000 3.075000 ;
      RECT 2.730000  0.085000 3.060000 0.700000 ;
      RECT 3.210000  1.875000 3.470000 2.735000 ;
      RECT 3.230000  0.255000 5.795000 0.425000 ;
      RECT 3.230000  0.425000 3.855000 0.870000 ;
      RECT 3.660000  2.035000 6.300000 2.205000 ;
      RECT 3.660000  2.205000 3.920000 2.905000 ;
      RECT 4.025000  0.595000 4.355000 0.870000 ;
      RECT 4.025000  0.870000 5.285000 1.040000 ;
      RECT 4.025000  1.040000 4.275000 1.185000 ;
      RECT 4.090000  2.375000 5.285000 2.545000 ;
      RECT 4.090000  2.545000 4.355000 3.075000 ;
      RECT 4.525000  0.425000 5.795000 0.435000 ;
      RECT 4.525000  0.435000 4.785000 0.700000 ;
      RECT 4.525000  2.715000 4.855000 3.245000 ;
      RECT 4.955000  0.615000 5.285000 0.870000 ;
      RECT 4.955000  1.040000 5.285000 1.075000 ;
      RECT 4.955000  1.075000 6.300000 1.255000 ;
      RECT 5.025000  2.545000 5.285000 3.075000 ;
      RECT 5.455000  2.205000 5.715000 3.075000 ;
      RECT 5.465000  0.435000 5.795000 0.895000 ;
      RECT 5.795000  1.255000 6.300000 1.395000 ;
      RECT 5.795000  1.395000 7.640000 1.585000 ;
      RECT 5.795000  1.585000 6.300000 2.035000 ;
      RECT 5.985000  0.085000 6.315000 0.905000 ;
      RECT 5.985000  2.375000 6.315000 3.245000 ;
      RECT 6.845000  0.085000 7.175000 0.885000 ;
      RECT 6.845000  2.095000 7.175000 3.245000 ;
      RECT 7.705000  0.085000 8.035000 0.885000 ;
      RECT 7.705000  2.095000 8.035000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_lp__o32a_4
END LIBRARY
