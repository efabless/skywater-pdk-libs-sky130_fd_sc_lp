# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__fa_0
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.504000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.870000 1.570000 2.950000 1.820000 ;
        RECT 0.870000 1.820000 1.120000 2.025000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.504000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.400000 1.990000 3.300000 2.320000 ;
        RECT 3.130000 1.755000 6.575000 1.925000 ;
        RECT 3.130000 1.925000 3.300000 1.990000 ;
        RECT 6.010000 1.925000 6.575000 2.125000 ;
        RECT 6.125000 1.190000 6.575000 1.755000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.690000 1.230000 3.790000 1.365000 ;
        RECT 1.690000 1.365000 5.835000 1.400000 ;
        RECT 3.435000 1.400000 5.835000 1.585000 ;
        RECT 3.450000 1.130000 3.790000 1.230000 ;
        RECT 5.505000 1.295000 5.835000 1.365000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.280900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.625000 0.495000 0.955000 ;
        RECT 0.085000 0.955000 0.325000 2.500000 ;
        RECT 0.085000 2.500000 0.425000 3.075000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.280900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.155000 0.350000 7.595000 0.680000 ;
        RECT 7.305000 1.405000 7.595000 2.945000 ;
        RECT 7.345000 0.680000 7.595000 1.405000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.495000  1.125000 1.520000 1.295000 ;
      RECT 0.495000  1.295000 0.700000 1.455000 ;
      RECT 0.530000  1.455000 0.700000 2.195000 ;
      RECT 0.530000  2.195000 1.230000 2.365000 ;
      RECT 0.595000  2.660000 0.890000 3.245000 ;
      RECT 0.665000  0.085000 0.995000 0.955000 ;
      RECT 1.060000  2.365000 1.230000 2.705000 ;
      RECT 1.060000  2.705000 1.825000 3.035000 ;
      RECT 1.255000  0.640000 1.745000 0.970000 ;
      RECT 1.255000  0.970000 1.520000 1.125000 ;
      RECT 1.915000  0.640000 2.245000 0.890000 ;
      RECT 1.915000  0.890000 3.235000 1.060000 ;
      RECT 1.995000  2.490000 3.225000 2.660000 ;
      RECT 1.995000  2.660000 2.275000 3.035000 ;
      RECT 2.415000  0.085000 2.745000 0.720000 ;
      RECT 2.445000  2.830000 2.775000 3.245000 ;
      RECT 2.915000  0.640000 3.235000 0.890000 ;
      RECT 2.945000  2.660000 3.225000 3.035000 ;
      RECT 3.450000  0.085000 3.780000 0.960000 ;
      RECT 3.470000  2.325000 3.745000 3.245000 ;
      RECT 3.915000  2.095000 5.145000 2.265000 ;
      RECT 3.915000  2.265000 4.190000 2.665000 ;
      RECT 3.960000  0.630000 4.190000 1.025000 ;
      RECT 3.960000  1.025000 5.140000 1.195000 ;
      RECT 4.360000  0.085000 4.690000 0.855000 ;
      RECT 4.360000  2.435000 4.690000 3.245000 ;
      RECT 4.860000  0.630000 5.140000 1.025000 ;
      RECT 4.860000  2.265000 5.145000 2.665000 ;
      RECT 5.310000  0.630000 5.600000 0.835000 ;
      RECT 5.310000  0.835000 6.520000 0.850000 ;
      RECT 5.310000  0.850000 7.175000 1.020000 ;
      RECT 5.315000  2.295000 6.955000 2.465000 ;
      RECT 5.315000  2.465000 5.645000 2.665000 ;
      RECT 6.690000  0.085000 6.985000 0.680000 ;
      RECT 6.745000  1.020000 7.175000 1.195000 ;
      RECT 6.745000  1.195000 6.955000 2.295000 ;
      RECT 6.805000  2.635000 7.135000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_lp__fa_0
END LIBRARY
