/*
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
*/


`ifndef SKY130_FD_SC_LP__O311AI_1_TIMING_V
`define SKY130_FD_SC_LP__O311AI_1_TIMING_V

/**
 * o311ai: 3-input OR into 3-input NAND.
 *
 *         Y = !((A1 | A2 | A3) & B1 & C1)
 *
 * Verilog simulation timing model.
 */

`timescale 1ns / 1ps
`default_nettype none

`celldefine
module sky130_fd_sc_lp__o311ai_1 (
    Y ,
    A1,
    A2,
    A3,
    B1,
    C1
);

    // Module ports
    output Y ;
    input  A1;
    input  A2;
    input  A3;
    input  B1;
    input  C1;

    // Module supplies
    supply1 VPWR;
    supply0 VGND;
    supply1 VPB ;
    supply0 VNB ;

    // Local signals
    wire or0_out    ;
    wire nand0_out_Y;

    //   Name   Output       Other arguments
    or   or0   (or0_out    , A2, A1, A3     );
    nand nand0 (nand0_out_Y, C1, or0_out, B1);
    buf  buf0  (Y          , nand0_out_Y    );

specify
(A1 -=> Y) = (0:0:0,0:0:0);
(A2 -=> Y) = (0:0:0,0:0:0);
(A3 -=> Y) = (0:0:0,0:0:0);
if ((!A1&!A2&A3&C1)) (B1 -=> Y) = (0:0:0,0:0:0);
if ((!A1&A2&!A3&C1)) (B1 -=> Y) = (0:0:0,0:0:0);
if ((!A1&A2&A3&C1)) (B1 -=> Y) = (0:0:0,0:0:0);
if ((A1&!A2&!A3&C1)) (B1 -=> Y) = (0:0:0,0:0:0);
if ((A1&!A2&A3&C1)) (B1 -=> Y) = (0:0:0,0:0:0);
if ((A1&A2&!A3&C1)) (B1 -=> Y) = (0:0:0,0:0:0);
if ((A1&A2&A3&C1)) (B1 -=> Y) = (0:0:0,0:0:0);
if ((!A1&!A2&A3&B1)) (C1 -=> Y) = (0:0:0,0:0:0);
if ((!A1&A2&!A3&B1)) (C1 -=> Y) = (0:0:0,0:0:0);
if ((!A1&A2&A3&B1)) (C1 -=> Y) = (0:0:0,0:0:0);
if ((A1&!A2&!A3&B1)) (C1 -=> Y) = (0:0:0,0:0:0);
if ((A1&!A2&A3&B1)) (C1 -=> Y) = (0:0:0,0:0:0);
if ((A1&A2&!A3&B1)) (C1 -=> Y) = (0:0:0,0:0:0);
if ((A1&A2&A3&B1)) (C1 -=> Y) = (0:0:0,0:0:0);
endspecify
endmodule
`endcelldefine

`default_nettype wire
`endif  // SKY130_FD_SC_LP__O311AI_1_TIMING_V
